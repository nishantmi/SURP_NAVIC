
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.CRFFT_pkg.ALL;

ENTITY TWDLROM IS
  PORT( clk                               :   IN    std_logic;
        reset                             :   IN    std_logic;
        enb                               :   IN    std_logic;
        dMemOutDly_vld                    :   IN    std_logic;
        stage                             :   IN    std_logic_vector(3 DOWNTO 0);  -- ufix4
        initIC                            :   IN    std_logic;
        syncReset                         :   IN    std_logic;
        twdl_re                           :   OUT   std_logic_vector(31 DOWNTO 0);  -- sfix32_En30
        twdl_im                           :   OUT   std_logic_vector(31 DOWNTO 0)  -- sfix32_En30
        );
END TWDLROM;


ARCHITECTURE rtl OF TWDLROM IS

  -- Constants
  CONSTANT Twiddle_re_table_data          : vector_of_signed32(0 TO 4095) := 
    (to_signed(1073741824, 32), to_signed(1073741804, 32), to_signed(1073741745, 32), to_signed(1073741646, 32),
     to_signed(1073741508, 32), to_signed(1073741331, 32), to_signed(1073741113, 32), to_signed(1073740857, 32),
     to_signed(1073740561, 32), to_signed(1073740225, 32), to_signed(1073739850, 32), to_signed(1073739436, 32),
     to_signed(1073738982, 32), to_signed(1073738488, 32), to_signed(1073737955, 32), to_signed(1073737383, 32),
     to_signed(1073736771, 32), to_signed(1073736119, 32), to_signed(1073735429, 32), to_signed(1073734698, 32),
     to_signed(1073733928, 32), to_signed(1073733119, 32), to_signed(1073732270, 32), to_signed(1073731382, 32),
     to_signed(1073730454, 32), to_signed(1073729487, 32), to_signed(1073728480, 32), to_signed(1073727434, 32),
     to_signed(1073726348, 32), to_signed(1073725223, 32), to_signed(1073724059, 32), to_signed(1073722855, 32),
     to_signed(1073721611, 32), to_signed(1073720328, 32), to_signed(1073719006, 32), to_signed(1073717644, 32),
     to_signed(1073716242, 32), to_signed(1073714801, 32), to_signed(1073713321, 32), to_signed(1073711801, 32),
     to_signed(1073710241, 32), to_signed(1073708643, 32), to_signed(1073707004, 32), to_signed(1073705326, 32),
     to_signed(1073703609, 32), to_signed(1073701852, 32), to_signed(1073700056, 32), to_signed(1073698220, 32),
     to_signed(1073696345, 32), to_signed(1073694431, 32), to_signed(1073692476, 32), to_signed(1073690483, 32),
     to_signed(1073688450, 32), to_signed(1073686377, 32), to_signed(1073684265, 32), to_signed(1073682113, 32),
     to_signed(1073679922, 32), to_signed(1073677692, 32), to_signed(1073675422, 32), to_signed(1073673113, 32),
     to_signed(1073670764, 32), to_signed(1073668375, 32), to_signed(1073665947, 32), to_signed(1073663480, 32),
     to_signed(1073660973, 32), to_signed(1073658427, 32), to_signed(1073655841, 32), to_signed(1073653216, 32),
     to_signed(1073650551, 32), to_signed(1073647847, 32), to_signed(1073645103, 32), to_signed(1073642320, 32),
     to_signed(1073639498, 32), to_signed(1073636635, 32), to_signed(1073633734, 32), to_signed(1073630793, 32),
     to_signed(1073627812, 32), to_signed(1073624792, 32), to_signed(1073621733, 32), to_signed(1073618634, 32),
     to_signed(1073615496, 32), to_signed(1073612318, 32), to_signed(1073609100, 32), to_signed(1073605843, 32),
     to_signed(1073602547, 32), to_signed(1073599211, 32), to_signed(1073595836, 32), to_signed(1073592421, 32),
     to_signed(1073588967, 32), to_signed(1073585474, 32), to_signed(1073581940, 32), to_signed(1073578368, 32),
     to_signed(1073574756, 32), to_signed(1073571104, 32), to_signed(1073567413, 32), to_signed(1073563683, 32),
     to_signed(1073559913, 32), to_signed(1073556103, 32), to_signed(1073552254, 32), to_signed(1073548366, 32),
     to_signed(1073544438, 32), to_signed(1073540471, 32), to_signed(1073536464, 32), to_signed(1073532418, 32),
     to_signed(1073528332, 32), to_signed(1073524207, 32), to_signed(1073520042, 32), to_signed(1073515838, 32),
     to_signed(1073511594, 32), to_signed(1073507311, 32), to_signed(1073502988, 32), to_signed(1073498626, 32),
     to_signed(1073494225, 32), to_signed(1073489784, 32), to_signed(1073485303, 32), to_signed(1073480784, 32),
     to_signed(1073476224, 32), to_signed(1073471625, 32), to_signed(1073466987, 32), to_signed(1073462309, 32),
     to_signed(1073457592, 32), to_signed(1073452835, 32), to_signed(1073448039, 32), to_signed(1073443203, 32),
     to_signed(1073438328, 32), to_signed(1073433414, 32), to_signed(1073428460, 32), to_signed(1073423466, 32),
     to_signed(1073418433, 32), to_signed(1073413361, 32), to_signed(1073408249, 32), to_signed(1073403097, 32),
     to_signed(1073397906, 32), to_signed(1073392676, 32), to_signed(1073387406, 32), to_signed(1073382097, 32),
     to_signed(1073376748, 32), to_signed(1073371360, 32), to_signed(1073365932, 32), to_signed(1073360465, 32),
     to_signed(1073354959, 32), to_signed(1073349413, 32), to_signed(1073343827, 32), to_signed(1073338202, 32),
     to_signed(1073332538, 32), to_signed(1073326834, 32), to_signed(1073321091, 32), to_signed(1073315308, 32),
     to_signed(1073309485, 32), to_signed(1073303624, 32), to_signed(1073297722, 32), to_signed(1073291782, 32),
     to_signed(1073285802, 32), to_signed(1073279782, 32), to_signed(1073273723, 32), to_signed(1073267624, 32),
     to_signed(1073261486, 32), to_signed(1073255309, 32), to_signed(1073249092, 32), to_signed(1073242836, 32),
     to_signed(1073236540, 32), to_signed(1073230205, 32), to_signed(1073223830, 32), to_signed(1073217416, 32),
     to_signed(1073210962, 32), to_signed(1073204469, 32), to_signed(1073197936, 32), to_signed(1073191364, 32),
     to_signed(1073184753, 32), to_signed(1073178102, 32), to_signed(1073171411, 32), to_signed(1073164682, 32),
     to_signed(1073157912, 32), to_signed(1073151103, 32), to_signed(1073144255, 32), to_signed(1073137367, 32),
     to_signed(1073130440, 32), to_signed(1073123474, 32), to_signed(1073116468, 32), to_signed(1073109422, 32),
     to_signed(1073102337, 32), to_signed(1073095213, 32), to_signed(1073088049, 32), to_signed(1073080845, 32),
     to_signed(1073073603, 32), to_signed(1073066320, 32), to_signed(1073058999, 32), to_signed(1073051638, 32),
     to_signed(1073044237, 32), to_signed(1073036797, 32), to_signed(1073029317, 32), to_signed(1073021798, 32),
     to_signed(1073014240, 32), to_signed(1073006642, 32), to_signed(1072999005, 32), to_signed(1072991328, 32),
     to_signed(1072983612, 32), to_signed(1072975856, 32), to_signed(1072968061, 32), to_signed(1072960226, 32),
     to_signed(1072952352, 32), to_signed(1072944439, 32), to_signed(1072936486, 32), to_signed(1072928494, 32),
     to_signed(1072920462, 32), to_signed(1072912391, 32), to_signed(1072904280, 32), to_signed(1072896130, 32),
     to_signed(1072887940, 32), to_signed(1072879711, 32), to_signed(1072871443, 32), to_signed(1072863135, 32),
     to_signed(1072854787, 32), to_signed(1072846400, 32), to_signed(1072837974, 32), to_signed(1072829508, 32),
     to_signed(1072821003, 32), to_signed(1072812458, 32), to_signed(1072803874, 32), to_signed(1072795251, 32),
     to_signed(1072786588, 32), to_signed(1072777886, 32), to_signed(1072769144, 32), to_signed(1072760362, 32),
     to_signed(1072751542, 32), to_signed(1072742682, 32), to_signed(1072733782, 32), to_signed(1072724843, 32),
     to_signed(1072715864, 32), to_signed(1072706846, 32), to_signed(1072697789, 32), to_signed(1072688692, 32),
     to_signed(1072679556, 32), to_signed(1072670380, 32), to_signed(1072661165, 32), to_signed(1072651911, 32),
     to_signed(1072642617, 32), to_signed(1072633283, 32), to_signed(1072623910, 32), to_signed(1072614498, 32),
     to_signed(1072605046, 32), to_signed(1072595555, 32), to_signed(1072586024, 32), to_signed(1072576454, 32),
     to_signed(1072566845, 32), to_signed(1072557196, 32), to_signed(1072547508, 32), to_signed(1072537780, 32),
     to_signed(1072528012, 32), to_signed(1072518206, 32), to_signed(1072508360, 32), to_signed(1072498474, 32),
     to_signed(1072488549, 32), to_signed(1072478585, 32), to_signed(1072468581, 32), to_signed(1072458538, 32),
     to_signed(1072448455, 32), to_signed(1072438333, 32), to_signed(1072428171, 32), to_signed(1072417970, 32),
     to_signed(1072407730, 32), to_signed(1072397450, 32), to_signed(1072387131, 32), to_signed(1072376772, 32),
     to_signed(1072366374, 32), to_signed(1072355936, 32), to_signed(1072345459, 32), to_signed(1072334943, 32),
     to_signed(1072324387, 32), to_signed(1072313792, 32), to_signed(1072303157, 32), to_signed(1072292483, 32),
     to_signed(1072281769, 32), to_signed(1072271016, 32), to_signed(1072260224, 32), to_signed(1072249392, 32),
     to_signed(1072238521, 32), to_signed(1072227610, 32), to_signed(1072216660, 32), to_signed(1072205671, 32),
     to_signed(1072194642, 32), to_signed(1072183573, 32), to_signed(1072172466, 32), to_signed(1072161318, 32),
     to_signed(1072150132, 32), to_signed(1072138906, 32), to_signed(1072127640, 32), to_signed(1072116335, 32),
     to_signed(1072104991, 32), to_signed(1072093607, 32), to_signed(1072082184, 32), to_signed(1072070722, 32),
     to_signed(1072059220, 32), to_signed(1072047678, 32), to_signed(1072036098, 32), to_signed(1072024477, 32),
     to_signed(1072012818, 32), to_signed(1072001119, 32), to_signed(1071989380, 32), to_signed(1071977602, 32),
     to_signed(1071965785, 32), to_signed(1071953928, 32), to_signed(1071942032, 32), to_signed(1071930097, 32),
     to_signed(1071918122, 32), to_signed(1071906107, 32), to_signed(1071894054, 32), to_signed(1071881960, 32),
     to_signed(1071869828, 32), to_signed(1071857656, 32), to_signed(1071845445, 32), to_signed(1071833194, 32),
     to_signed(1071820903, 32), to_signed(1071808574, 32), to_signed(1071796205, 32), to_signed(1071783796, 32),
     to_signed(1071771349, 32), to_signed(1071758861, 32), to_signed(1071746335, 32), to_signed(1071733769, 32),
     to_signed(1071721163, 32), to_signed(1071708518, 32), to_signed(1071695834, 32), to_signed(1071683110, 32),
     to_signed(1071670347, 32), to_signed(1071657545, 32), to_signed(1071644703, 32), to_signed(1071631822, 32),
     to_signed(1071618901, 32), to_signed(1071605941, 32), to_signed(1071592941, 32), to_signed(1071579902, 32),
     to_signed(1071566824, 32), to_signed(1071553706, 32), to_signed(1071540549, 32), to_signed(1071527353, 32),
     to_signed(1071514117, 32), to_signed(1071500842, 32), to_signed(1071487527, 32), to_signed(1071474173, 32),
     to_signed(1071460780, 32), to_signed(1071447347, 32), to_signed(1071433874, 32), to_signed(1071420363, 32),
     to_signed(1071406812, 32), to_signed(1071393221, 32), to_signed(1071379592, 32), to_signed(1071365922, 32),
     to_signed(1071352214, 32), to_signed(1071338466, 32), to_signed(1071324678, 32), to_signed(1071310852, 32),
     to_signed(1071296985, 32), to_signed(1071283080, 32), to_signed(1071269135, 32), to_signed(1071255151, 32),
     to_signed(1071241127, 32), to_signed(1071227064, 32), to_signed(1071212961, 32), to_signed(1071198819, 32),
     to_signed(1071184638, 32), to_signed(1071170418, 32), to_signed(1071156158, 32), to_signed(1071141858, 32),
     to_signed(1071127519, 32), to_signed(1071113141, 32), to_signed(1071098724, 32), to_signed(1071084267, 32),
     to_signed(1071069770, 32), to_signed(1071055235, 32), to_signed(1071040660, 32), to_signed(1071026045, 32),
     to_signed(1071011391, 32), to_signed(1070996698, 32), to_signed(1070981966, 32), to_signed(1070967194, 32),
     to_signed(1070952382, 32), to_signed(1070937532, 32), to_signed(1070922641, 32), to_signed(1070907712, 32),
     to_signed(1070892743, 32), to_signed(1070877735, 32), to_signed(1070862687, 32), to_signed(1070847600, 32),
     to_signed(1070832474, 32), to_signed(1070817308, 32), to_signed(1070802103, 32), to_signed(1070786859, 32),
     to_signed(1070771575, 32), to_signed(1070756252, 32), to_signed(1070740889, 32), to_signed(1070725487, 32),
     to_signed(1070710046, 32), to_signed(1070694565, 32), to_signed(1070679045, 32), to_signed(1070663486, 32),
     to_signed(1070647887, 32), to_signed(1070632249, 32), to_signed(1070616572, 32), to_signed(1070600855, 32),
     to_signed(1070585099, 32), to_signed(1070569303, 32), to_signed(1070553468, 32), to_signed(1070537594, 32),
     to_signed(1070521680, 32), to_signed(1070505727, 32), to_signed(1070489735, 32), to_signed(1070473703, 32),
     to_signed(1070457632, 32), to_signed(1070441521, 32), to_signed(1070425372, 32), to_signed(1070409182, 32),
     to_signed(1070392954, 32), to_signed(1070376686, 32), to_signed(1070360379, 32), to_signed(1070344032, 32),
     to_signed(1070327646, 32), to_signed(1070311221, 32), to_signed(1070294756, 32), to_signed(1070278252, 32),
     to_signed(1070261709, 32), to_signed(1070245126, 32), to_signed(1070228504, 32), to_signed(1070211843, 32),
     to_signed(1070195142, 32), to_signed(1070178402, 32), to_signed(1070161623, 32), to_signed(1070144804, 32),
     to_signed(1070127946, 32), to_signed(1070111048, 32), to_signed(1070094111, 32), to_signed(1070077135, 32),
     to_signed(1070060120, 32), to_signed(1070043065, 32), to_signed(1070025971, 32), to_signed(1070008837, 32),
     to_signed(1069991664, 32), to_signed(1069974452, 32), to_signed(1069957201, 32), to_signed(1069939910, 32),
     to_signed(1069922579, 32), to_signed(1069905210, 32), to_signed(1069887801, 32), to_signed(1069870353, 32),
     to_signed(1069852865, 32), to_signed(1069835338, 32), to_signed(1069817772, 32), to_signed(1069800166, 32),
     to_signed(1069782521, 32), to_signed(1069764837, 32), to_signed(1069747114, 32), to_signed(1069729351, 32),
     to_signed(1069711548, 32), to_signed(1069693707, 32), to_signed(1069675826, 32), to_signed(1069657906, 32),
     to_signed(1069639946, 32), to_signed(1069621947, 32), to_signed(1069603909, 32), to_signed(1069585832, 32),
     to_signed(1069567715, 32), to_signed(1069549558, 32), to_signed(1069531363, 32), to_signed(1069513128, 32),
     to_signed(1069494854, 32), to_signed(1069476540, 32), to_signed(1069458188, 32), to_signed(1069439795, 32),
     to_signed(1069421364, 32), to_signed(1069402893, 32), to_signed(1069384383, 32), to_signed(1069365834, 32),
     to_signed(1069347245, 32), to_signed(1069328617, 32), to_signed(1069309950, 32), to_signed(1069291243, 32),
     to_signed(1069272497, 32), to_signed(1069253712, 32), to_signed(1069234887, 32), to_signed(1069216023, 32),
     to_signed(1069197120, 32), to_signed(1069178177, 32), to_signed(1069159195, 32), to_signed(1069140174, 32),
     to_signed(1069121114, 32), to_signed(1069102014, 32), to_signed(1069082875, 32), to_signed(1069063697, 32),
     to_signed(1069044479, 32), to_signed(1069025222, 32), to_signed(1069005925, 32), to_signed(1068986590, 32),
     to_signed(1068967215, 32), to_signed(1068947801, 32), to_signed(1068928347, 32), to_signed(1068908854, 32),
     to_signed(1068889322, 32), to_signed(1068869751, 32), to_signed(1068850140, 32), to_signed(1068830490, 32),
     to_signed(1068810801, 32), to_signed(1068791072, 32), to_signed(1068771304, 32), to_signed(1068751497, 32),
     to_signed(1068731650, 32), to_signed(1068711764, 32), to_signed(1068691839, 32), to_signed(1068671875, 32),
     to_signed(1068651871, 32), to_signed(1068631828, 32), to_signed(1068611746, 32), to_signed(1068591624, 32),
     to_signed(1068571464, 32), to_signed(1068551263, 32), to_signed(1068531024, 32), to_signed(1068510745, 32),
     to_signed(1068490427, 32), to_signed(1068470070, 32), to_signed(1068449673, 32), to_signed(1068429238, 32),
     to_signed(1068408763, 32), to_signed(1068388248, 32), to_signed(1068367694, 32), to_signed(1068347101, 32),
     to_signed(1068326469, 32), to_signed(1068305798, 32), to_signed(1068285087, 32), to_signed(1068264337, 32),
     to_signed(1068243547, 32), to_signed(1068222719, 32), to_signed(1068201851, 32), to_signed(1068180944, 32),
     to_signed(1068159997, 32), to_signed(1068139011, 32), to_signed(1068117986, 32), to_signed(1068096922, 32),
     to_signed(1068075818, 32), to_signed(1068054676, 32), to_signed(1068033493, 32), to_signed(1068012272, 32),
     to_signed(1067991011, 32), to_signed(1067969712, 32), to_signed(1067948372, 32), to_signed(1067926994, 32),
     to_signed(1067905576, 32), to_signed(1067884119, 32), to_signed(1067862623, 32), to_signed(1067841088, 32),
     to_signed(1067819513, 32), to_signed(1067797899, 32), to_signed(1067776246, 32), to_signed(1067754553, 32),
     to_signed(1067732821, 32), to_signed(1067711050, 32), to_signed(1067689240, 32), to_signed(1067667390, 32),
     to_signed(1067645501, 32), to_signed(1067623573, 32), to_signed(1067601606, 32), to_signed(1067579600, 32),
     to_signed(1067557554, 32), to_signed(1067535469, 32), to_signed(1067513344, 32), to_signed(1067491181, 32),
     to_signed(1067468978, 32), to_signed(1067446736, 32), to_signed(1067424454, 32), to_signed(1067402134, 32),
     to_signed(1067379774, 32), to_signed(1067357375, 32), to_signed(1067334937, 32), to_signed(1067312459, 32),
     to_signed(1067289942, 32), to_signed(1067267386, 32), to_signed(1067244791, 32), to_signed(1067222157, 32),
     to_signed(1067199483, 32), to_signed(1067176770, 32), to_signed(1067154018, 32), to_signed(1067131226, 32),
     to_signed(1067108396, 32), to_signed(1067085526, 32), to_signed(1067062616, 32), to_signed(1067039668, 32),
     to_signed(1067016680, 32), to_signed(1066993654, 32), to_signed(1066970587, 32), to_signed(1066947482, 32),
     to_signed(1066924338, 32), to_signed(1066901154, 32), to_signed(1066877931, 32), to_signed(1066854669, 32),
     to_signed(1066831367, 32), to_signed(1066808026, 32), to_signed(1066784647, 32), to_signed(1066761227, 32),
     to_signed(1066737769, 32), to_signed(1066714272, 32), to_signed(1066690735, 32), to_signed(1066667159, 32),
     to_signed(1066643544, 32), to_signed(1066619889, 32), to_signed(1066596195, 32), to_signed(1066572463, 32),
     to_signed(1066548690, 32), to_signed(1066524879, 32), to_signed(1066501029, 32), to_signed(1066477139, 32),
     to_signed(1066453210, 32), to_signed(1066429242, 32), to_signed(1066405234, 32), to_signed(1066381188, 32),
     to_signed(1066357102, 32), to_signed(1066332977, 32), to_signed(1066308813, 32), to_signed(1066284610, 32),
     to_signed(1066260367, 32), to_signed(1066236085, 32), to_signed(1066211764, 32), to_signed(1066187404, 32),
     to_signed(1066163005, 32), to_signed(1066138566, 32), to_signed(1066114088, 32), to_signed(1066089571, 32),
     to_signed(1066065015, 32), to_signed(1066040420, 32), to_signed(1066015785, 32), to_signed(1065991111, 32),
     to_signed(1065966398, 32), to_signed(1065941646, 32), to_signed(1065916855, 32), to_signed(1065892024, 32),
     to_signed(1065867154, 32), to_signed(1065842245, 32), to_signed(1065817297, 32), to_signed(1065792310, 32),
     to_signed(1065767284, 32), to_signed(1065742218, 32), to_signed(1065717113, 32), to_signed(1065691969, 32),
     to_signed(1065666786, 32), to_signed(1065641563, 32), to_signed(1065616302, 32), to_signed(1065591001, 32),
     to_signed(1065565661, 32), to_signed(1065540282, 32), to_signed(1065514864, 32), to_signed(1065489406, 32),
     to_signed(1065463909, 32), to_signed(1065438374, 32), to_signed(1065412799, 32), to_signed(1065387184, 32),
     to_signed(1065361531, 32), to_signed(1065335839, 32), to_signed(1065310107, 32), to_signed(1065284336, 32),
     to_signed(1065258526, 32), to_signed(1065232677, 32), to_signed(1065206789, 32), to_signed(1065180861, 32),
     to_signed(1065154894, 32), to_signed(1065128889, 32), to_signed(1065102844, 32), to_signed(1065076759, 32),
     to_signed(1065050636, 32), to_signed(1065024474, 32), to_signed(1064998272, 32), to_signed(1064972031, 32),
     to_signed(1064945751, 32), to_signed(1064919432, 32), to_signed(1064893074, 32), to_signed(1064866676, 32),
     to_signed(1064840240, 32), to_signed(1064813764, 32), to_signed(1064787249, 32), to_signed(1064760695, 32),
     to_signed(1064734102, 32), to_signed(1064707470, 32), to_signed(1064680798, 32), to_signed(1064654088, 32),
     to_signed(1064627338, 32), to_signed(1064600549, 32), to_signed(1064573721, 32), to_signed(1064546854, 32),
     to_signed(1064519947, 32), to_signed(1064493002, 32), to_signed(1064466017, 32), to_signed(1064438994, 32),
     to_signed(1064411931, 32), to_signed(1064384829, 32), to_signed(1064357688, 32), to_signed(1064330507, 32),
     to_signed(1064303288, 32), to_signed(1064276029, 32), to_signed(1064248732, 32), to_signed(1064221395, 32),
     to_signed(1064194019, 32), to_signed(1064166604, 32), to_signed(1064139150, 32), to_signed(1064111657, 32),
     to_signed(1064084124, 32), to_signed(1064056553, 32), to_signed(1064028942, 32), to_signed(1064001292, 32),
     to_signed(1063973603, 32), to_signed(1063945875, 32), to_signed(1063918108, 32), to_signed(1063890302, 32),
     to_signed(1063862456, 32), to_signed(1063834572, 32), to_signed(1063806648, 32), to_signed(1063778685, 32),
     to_signed(1063750684, 32), to_signed(1063722643, 32), to_signed(1063694563, 32), to_signed(1063666443, 32),
     to_signed(1063638285, 32), to_signed(1063610088, 32), to_signed(1063581851, 32), to_signed(1063553576, 32),
     to_signed(1063525261, 32), to_signed(1063496907, 32), to_signed(1063468514, 32), to_signed(1063440082, 32),
     to_signed(1063411611, 32), to_signed(1063383101, 32), to_signed(1063354552, 32), to_signed(1063325963, 32),
     to_signed(1063297336, 32), to_signed(1063268669, 32), to_signed(1063239964, 32), to_signed(1063211219, 32),
     to_signed(1063182435, 32), to_signed(1063153612, 32), to_signed(1063124750, 32), to_signed(1063095849, 32),
     to_signed(1063066909, 32), to_signed(1063037929, 32), to_signed(1063008911, 32), to_signed(1062979853, 32),
     to_signed(1062950757, 32), to_signed(1062921621, 32), to_signed(1062892446, 32), to_signed(1062863233, 32),
     to_signed(1062833980, 32), to_signed(1062804688, 32), to_signed(1062775357, 32), to_signed(1062745987, 32),
     to_signed(1062716578, 32), to_signed(1062687129, 32), to_signed(1062657642, 32), to_signed(1062628116, 32),
     to_signed(1062598550, 32), to_signed(1062568946, 32), to_signed(1062539302, 32), to_signed(1062509619, 32),
     to_signed(1062479898, 32), to_signed(1062450137, 32), to_signed(1062420337, 32), to_signed(1062390498, 32),
     to_signed(1062360620, 32), to_signed(1062330703, 32), to_signed(1062300747, 32), to_signed(1062270752, 32),
     to_signed(1062240717, 32), to_signed(1062210644, 32), to_signed(1062180532, 32), to_signed(1062150381, 32),
     to_signed(1062120190, 32), to_signed(1062089961, 32), to_signed(1062059692, 32), to_signed(1062029384, 32),
     to_signed(1061999038, 32), to_signed(1061968652, 32), to_signed(1061938227, 32), to_signed(1061907764, 32),
     to_signed(1061877261, 32), to_signed(1061846719, 32), to_signed(1061816138, 32), to_signed(1061785518, 32),
     to_signed(1061754859, 32), to_signed(1061724161, 32), to_signed(1061693424, 32), to_signed(1061662648, 32),
     to_signed(1061631833, 32), to_signed(1061600979, 32), to_signed(1061570086, 32), to_signed(1061539153, 32),
     to_signed(1061508182, 32), to_signed(1061477172, 32), to_signed(1061446123, 32), to_signed(1061415034, 32),
     to_signed(1061383907, 32), to_signed(1061352741, 32), to_signed(1061321535, 32), to_signed(1061290291, 32),
     to_signed(1061259007, 32), to_signed(1061227685, 32), to_signed(1061196323, 32), to_signed(1061164923, 32),
     to_signed(1061133483, 32), to_signed(1061102005, 32), to_signed(1061070487, 32), to_signed(1061038931, 32),
     to_signed(1061007335, 32), to_signed(1060975701, 32), to_signed(1060944027, 32), to_signed(1060912314, 32),
     to_signed(1060880563, 32), to_signed(1060848772, 32), to_signed(1060816943, 32), to_signed(1060785074, 32),
     to_signed(1060753166, 32), to_signed(1060721220, 32), to_signed(1060689234, 32), to_signed(1060657210, 32),
     to_signed(1060625146, 32), to_signed(1060593043, 32), to_signed(1060560902, 32), to_signed(1060528721, 32),
     to_signed(1060496502, 32), to_signed(1060464243, 32), to_signed(1060431945, 32), to_signed(1060399609, 32),
     to_signed(1060367233, 32), to_signed(1060334819, 32), to_signed(1060302365, 32), to_signed(1060269873, 32),
     to_signed(1060237341, 32), to_signed(1060204771, 32), to_signed(1060172161, 32), to_signed(1060139513, 32),
     to_signed(1060106826, 32), to_signed(1060074099, 32), to_signed(1060041334, 32), to_signed(1060008530, 32),
     to_signed(1059975686, 32), to_signed(1059942804, 32), to_signed(1059909883, 32), to_signed(1059876922, 32),
     to_signed(1059843923, 32), to_signed(1059810885, 32), to_signed(1059777808, 32), to_signed(1059744692, 32),
     to_signed(1059711537, 32), to_signed(1059678343, 32), to_signed(1059645110, 32), to_signed(1059611838, 32),
     to_signed(1059578527, 32), to_signed(1059545177, 32), to_signed(1059511788, 32), to_signed(1059478361, 32),
     to_signed(1059444894, 32), to_signed(1059411388, 32), to_signed(1059377844, 32), to_signed(1059344260, 32),
     to_signed(1059310638, 32), to_signed(1059276976, 32), to_signed(1059243276, 32), to_signed(1059209536, 32),
     to_signed(1059175758, 32), to_signed(1059141941, 32), to_signed(1059108085, 32), to_signed(1059074189, 32),
     to_signed(1059040255, 32), to_signed(1059006282, 32), to_signed(1058972270, 32), to_signed(1058938220, 32),
     to_signed(1058904130, 32), to_signed(1058870001, 32), to_signed(1058835833, 32), to_signed(1058801627, 32),
     to_signed(1058767381, 32), to_signed(1058733097, 32), to_signed(1058698773, 32), to_signed(1058664411, 32),
     to_signed(1058630010, 32), to_signed(1058595570, 32), to_signed(1058561091, 32), to_signed(1058526573, 32),
     to_signed(1058492016, 32), to_signed(1058457420, 32), to_signed(1058422785, 32), to_signed(1058388111, 32),
     to_signed(1058353399, 32), to_signed(1058318647, 32), to_signed(1058283857, 32), to_signed(1058249028, 32),
     to_signed(1058214159, 32), to_signed(1058179252, 32), to_signed(1058144306, 32), to_signed(1058109321, 32),
     to_signed(1058074297, 32), to_signed(1058039235, 32), to_signed(1058004133, 32), to_signed(1057968992, 32),
     to_signed(1057933813, 32), to_signed(1057898595, 32), to_signed(1057863337, 32), to_signed(1057828041, 32),
     to_signed(1057792706, 32), to_signed(1057757332, 32), to_signed(1057721919, 32), to_signed(1057686468, 32),
     to_signed(1057650977, 32), to_signed(1057615448, 32), to_signed(1057579879, 32), to_signed(1057544272, 32),
     to_signed(1057508626, 32), to_signed(1057472941, 32), to_signed(1057437217, 32), to_signed(1057401454, 32),
     to_signed(1057365653, 32), to_signed(1057329812, 32), to_signed(1057293933, 32), to_signed(1057258014, 32),
     to_signed(1057222057, 32), to_signed(1057186061, 32), to_signed(1057150026, 32), to_signed(1057113952, 32),
     to_signed(1057077840, 32), to_signed(1057041688, 32), to_signed(1057005498, 32), to_signed(1056969269, 32),
     to_signed(1056933001, 32), to_signed(1056896694, 32), to_signed(1056860348, 32), to_signed(1056823963, 32),
     to_signed(1056787540, 32), to_signed(1056751077, 32), to_signed(1056714576, 32), to_signed(1056678036, 32),
     to_signed(1056641457, 32), to_signed(1056604839, 32), to_signed(1056568183, 32), to_signed(1056531487, 32),
     to_signed(1056494753, 32), to_signed(1056457980, 32), to_signed(1056421168, 32), to_signed(1056384317, 32),
     to_signed(1056347427, 32), to_signed(1056310499, 32), to_signed(1056273531, 32), to_signed(1056236525, 32),
     to_signed(1056199480, 32), to_signed(1056162396, 32), to_signed(1056125274, 32), to_signed(1056088112, 32),
     to_signed(1056050912, 32), to_signed(1056013673, 32), to_signed(1055976395, 32), to_signed(1055939078, 32),
     to_signed(1055901722, 32), to_signed(1055864328, 32), to_signed(1055826894, 32), to_signed(1055789422, 32),
     to_signed(1055751911, 32), to_signed(1055714361, 32), to_signed(1055676773, 32), to_signed(1055639145, 32),
     to_signed(1055601479, 32), to_signed(1055563774, 32), to_signed(1055526030, 32), to_signed(1055488248, 32),
     to_signed(1055450426, 32), to_signed(1055412566, 32), to_signed(1055374667, 32), to_signed(1055336729, 32),
     to_signed(1055298753, 32), to_signed(1055260737, 32), to_signed(1055222683, 32), to_signed(1055184590, 32),
     to_signed(1055146458, 32), to_signed(1055108287, 32), to_signed(1055070078, 32), to_signed(1055031830, 32),
     to_signed(1054993543, 32), to_signed(1054955217, 32), to_signed(1054916852, 32), to_signed(1054878449, 32),
     to_signed(1054840007, 32), to_signed(1054801526, 32), to_signed(1054763006, 32), to_signed(1054724447, 32),
     to_signed(1054685850, 32), to_signed(1054647214, 32), to_signed(1054608539, 32), to_signed(1054569826, 32),
     to_signed(1054531073, 32), to_signed(1054492282, 32), to_signed(1054453452, 32), to_signed(1054414583, 32),
     to_signed(1054375676, 32), to_signed(1054336730, 32), to_signed(1054297745, 32), to_signed(1054258721, 32),
     to_signed(1054219658, 32), to_signed(1054180557, 32), to_signed(1054141417, 32), to_signed(1054102238, 32),
     to_signed(1054063021, 32), to_signed(1054023764, 32), to_signed(1053984469, 32), to_signed(1053945135, 32),
     to_signed(1053905763, 32), to_signed(1053866352, 32), to_signed(1053826901, 32), to_signed(1053787413, 32),
     to_signed(1053747885, 32), to_signed(1053708319, 32), to_signed(1053668714, 32), to_signed(1053629070, 32),
     to_signed(1053589387, 32), to_signed(1053549666, 32), to_signed(1053509906, 32), to_signed(1053470107, 32),
     to_signed(1053430270, 32), to_signed(1053390394, 32), to_signed(1053350479, 32), to_signed(1053310525, 32),
     to_signed(1053270533, 32), to_signed(1053230502, 32), to_signed(1053190432, 32), to_signed(1053150323, 32),
     to_signed(1053110176, 32), to_signed(1053069990, 32), to_signed(1053029765, 32), to_signed(1052989502, 32),
     to_signed(1052949200, 32), to_signed(1052908859, 32), to_signed(1052868479, 32), to_signed(1052828061, 32),
     to_signed(1052787604, 32), to_signed(1052747108, 32), to_signed(1052706574, 32), to_signed(1052666001, 32),
     to_signed(1052625389, 32), to_signed(1052584738, 32), to_signed(1052544049, 32), to_signed(1052503321, 32),
     to_signed(1052462555, 32), to_signed(1052421749, 32), to_signed(1052380905, 32), to_signed(1052340022, 32),
     to_signed(1052299101, 32), to_signed(1052258141, 32), to_signed(1052217142, 32), to_signed(1052176105, 32),
     to_signed(1052135029, 32), to_signed(1052093914, 32), to_signed(1052052760, 32), to_signed(1052011568, 32),
     to_signed(1051970337, 32), to_signed(1051929068, 32), to_signed(1051887759, 32), to_signed(1051846413, 32),
     to_signed(1051805027, 32), to_signed(1051763603, 32), to_signed(1051722140, 32), to_signed(1051680638, 32),
     to_signed(1051639098, 32), to_signed(1051597519, 32), to_signed(1051555901, 32), to_signed(1051514245, 32),
     to_signed(1051472550, 32), to_signed(1051430817, 32), to_signed(1051389044, 32), to_signed(1051347234, 32),
     to_signed(1051305384, 32), to_signed(1051263496, 32), to_signed(1051221569, 32), to_signed(1051179604, 32),
     to_signed(1051137599, 32), to_signed(1051095557, 32), to_signed(1051053475, 32), to_signed(1051011355, 32),
     to_signed(1050969196, 32), to_signed(1050926999, 32), to_signed(1050884763, 32), to_signed(1050842488, 32),
     to_signed(1050800175, 32), to_signed(1050757823, 32), to_signed(1050715433, 32), to_signed(1050673003, 32),
     to_signed(1050630536, 32), to_signed(1050588029, 32), to_signed(1050545484, 32), to_signed(1050502900, 32),
     to_signed(1050460278, 32), to_signed(1050417617, 32), to_signed(1050374918, 32), to_signed(1050332179, 32),
     to_signed(1050289403, 32), to_signed(1050246587, 32), to_signed(1050203733, 32), to_signed(1050160841, 32),
     to_signed(1050117909, 32), to_signed(1050074939, 32), to_signed(1050031931, 32), to_signed(1049988884, 32),
     to_signed(1049945798, 32), to_signed(1049902674, 32), to_signed(1049859511, 32), to_signed(1049816310, 32),
     to_signed(1049773069, 32), to_signed(1049729791, 32), to_signed(1049686474, 32), to_signed(1049643118, 32),
     to_signed(1049599723, 32), to_signed(1049556290, 32), to_signed(1049512818, 32), to_signed(1049469308, 32),
     to_signed(1049425759, 32), to_signed(1049382172, 32), to_signed(1049338546, 32), to_signed(1049294881, 32),
     to_signed(1049251178, 32), to_signed(1049207437, 32), to_signed(1049163656, 32), to_signed(1049119837, 32),
     to_signed(1049075980, 32), to_signed(1049032084, 32), to_signed(1048988149, 32), to_signed(1048944176, 32),
     to_signed(1048900165, 32), to_signed(1048856114, 32), to_signed(1048812025, 32), to_signed(1048767898, 32),
     to_signed(1048723732, 32), to_signed(1048679527, 32), to_signed(1048635284, 32), to_signed(1048591003, 32),
     to_signed(1048546683, 32), to_signed(1048502324, 32), to_signed(1048457926, 32), to_signed(1048413491, 32),
     to_signed(1048369016, 32), to_signed(1048324503, 32), to_signed(1048279952, 32), to_signed(1048235362, 32),
     to_signed(1048190733, 32), to_signed(1048146066, 32), to_signed(1048101360, 32), to_signed(1048056616, 32),
     to_signed(1048011834, 32), to_signed(1047967012, 32), to_signed(1047922153, 32), to_signed(1047877254, 32),
     to_signed(1047832317, 32), to_signed(1047787342, 32), to_signed(1047742328, 32), to_signed(1047697276, 32),
     to_signed(1047652185, 32), to_signed(1047607055, 32), to_signed(1047561887, 32), to_signed(1047516681, 32),
     to_signed(1047471436, 32), to_signed(1047426152, 32), to_signed(1047380830, 32), to_signed(1047335470, 32),
     to_signed(1047290071, 32), to_signed(1047244633, 32), to_signed(1047199157, 32), to_signed(1047153643, 32),
     to_signed(1047108090, 32), to_signed(1047062498, 32), to_signed(1047016868, 32), to_signed(1046971199, 32),
     to_signed(1046925492, 32), to_signed(1046879747, 32), to_signed(1046833963, 32), to_signed(1046788140, 32),
     to_signed(1046742279, 32), to_signed(1046696380, 32), to_signed(1046650442, 32), to_signed(1046604466, 32),
     to_signed(1046558451, 32), to_signed(1046512397, 32), to_signed(1046466305, 32), to_signed(1046420175, 32),
     to_signed(1046374006, 32), to_signed(1046327799, 32), to_signed(1046281553, 32), to_signed(1046235269, 32),
     to_signed(1046188946, 32), to_signed(1046142585, 32), to_signed(1046096185, 32), to_signed(1046049747, 32),
     to_signed(1046003271, 32), to_signed(1045956756, 32), to_signed(1045910202, 32), to_signed(1045863610, 32),
     to_signed(1045816980, 32), to_signed(1045770311, 32), to_signed(1045723604, 32), to_signed(1045676858, 32),
     to_signed(1045630074, 32), to_signed(1045583251, 32), to_signed(1045536390, 32), to_signed(1045489490, 32),
     to_signed(1045442553, 32), to_signed(1045395576, 32), to_signed(1045348561, 32), to_signed(1045301508, 32),
     to_signed(1045254416, 32), to_signed(1045207286, 32), to_signed(1045160118, 32), to_signed(1045112911, 32),
     to_signed(1045065665, 32), to_signed(1045018381, 32), to_signed(1044971059, 32), to_signed(1044923699, 32),
     to_signed(1044876299, 32), to_signed(1044828862, 32), to_signed(1044781386, 32), to_signed(1044733872, 32),
     to_signed(1044686319, 32), to_signed(1044638728, 32), to_signed(1044591098, 32), to_signed(1044543430, 32),
     to_signed(1044495724, 32), to_signed(1044447979, 32), to_signed(1044400196, 32), to_signed(1044352374, 32),
     to_signed(1044304514, 32), to_signed(1044256616, 32), to_signed(1044208679, 32), to_signed(1044160704, 32),
     to_signed(1044112690, 32), to_signed(1044064638, 32), to_signed(1044016548, 32), to_signed(1043968419, 32),
     to_signed(1043920252, 32), to_signed(1043872047, 32), to_signed(1043823803, 32), to_signed(1043775521, 32),
     to_signed(1043727200, 32), to_signed(1043678841, 32), to_signed(1043630444, 32), to_signed(1043582008, 32),
     to_signed(1043533534, 32), to_signed(1043485021, 32), to_signed(1043436471, 32), to_signed(1043387881, 32),
     to_signed(1043339254, 32), to_signed(1043290588, 32), to_signed(1043241884, 32), to_signed(1043193141, 32),
     to_signed(1043144360, 32), to_signed(1043095541, 32), to_signed(1043046683, 32), to_signed(1042997787, 32),
     to_signed(1042948852, 32), to_signed(1042899880, 32), to_signed(1042850869, 32), to_signed(1042801819, 32),
     to_signed(1042752731, 32), to_signed(1042703605, 32), to_signed(1042654441, 32), to_signed(1042605238, 32),
     to_signed(1042555997, 32), to_signed(1042506717, 32), to_signed(1042457400, 32), to_signed(1042408044, 32),
     to_signed(1042358649, 32), to_signed(1042309216, 32), to_signed(1042259745, 32), to_signed(1042210236, 32),
     to_signed(1042160688, 32), to_signed(1042111102, 32), to_signed(1042061478, 32), to_signed(1042011815, 32),
     to_signed(1041962114, 32), to_signed(1041912375, 32), to_signed(1041862597, 32), to_signed(1041812781, 32),
     to_signed(1041762927, 32), to_signed(1041713034, 32), to_signed(1041663104, 32), to_signed(1041613135, 32),
     to_signed(1041563127, 32), to_signed(1041513081, 32), to_signed(1041462997, 32), to_signed(1041412875, 32),
     to_signed(1041362715, 32), to_signed(1041312516, 32), to_signed(1041262279, 32), to_signed(1041212003, 32),
     to_signed(1041161689, 32), to_signed(1041111337, 32), to_signed(1041060947, 32), to_signed(1041010519, 32),
     to_signed(1040960052, 32), to_signed(1040909547, 32), to_signed(1040859003, 32), to_signed(1040808422, 32),
     to_signed(1040757802, 32), to_signed(1040707143, 32), to_signed(1040656447, 32), to_signed(1040605712, 32),
     to_signed(1040554939, 32), to_signed(1040504128, 32), to_signed(1040453279, 32), to_signed(1040402391, 32),
     to_signed(1040351465, 32), to_signed(1040300501, 32), to_signed(1040249498, 32), to_signed(1040198457, 32),
     to_signed(1040147378, 32), to_signed(1040096261, 32), to_signed(1040045106, 32), to_signed(1039993912, 32),
     to_signed(1039942680, 32), to_signed(1039891410, 32), to_signed(1039840101, 32), to_signed(1039788755, 32),
     to_signed(1039737370, 32), to_signed(1039685947, 32), to_signed(1039634486, 32), to_signed(1039582986, 32),
     to_signed(1039531448, 32), to_signed(1039479872, 32), to_signed(1039428258, 32), to_signed(1039376606, 32),
     to_signed(1039324915, 32), to_signed(1039273186, 32), to_signed(1039221419, 32), to_signed(1039169614, 32),
     to_signed(1039117770, 32), to_signed(1039065889, 32), to_signed(1039013969, 32), to_signed(1038962011, 32),
     to_signed(1038910014, 32), to_signed(1038857980, 32), to_signed(1038805907, 32), to_signed(1038753796, 32),
     to_signed(1038701647, 32), to_signed(1038649460, 32), to_signed(1038597234, 32), to_signed(1038544971, 32),
     to_signed(1038492669, 32), to_signed(1038440329, 32), to_signed(1038387951, 32), to_signed(1038335534, 32),
     to_signed(1038283080, 32), to_signed(1038230587, 32), to_signed(1038178056, 32), to_signed(1038125487, 32),
     to_signed(1038072880, 32), to_signed(1038020234, 32), to_signed(1037967551, 32), to_signed(1037914829, 32),
     to_signed(1037862069, 32), to_signed(1037809271, 32), to_signed(1037756435, 32), to_signed(1037703561, 32),
     to_signed(1037650648, 32), to_signed(1037597698, 32), to_signed(1037544709, 32), to_signed(1037491682, 32),
     to_signed(1037438617, 32), to_signed(1037385513, 32), to_signed(1037332372, 32), to_signed(1037279192, 32),
     to_signed(1037225975, 32), to_signed(1037172719, 32), to_signed(1037119425, 32), to_signed(1037066093, 32),
     to_signed(1037012723, 32), to_signed(1036959314, 32), to_signed(1036905868, 32), to_signed(1036852383, 32),
     to_signed(1036798861, 32), to_signed(1036745300, 32), to_signed(1036691701, 32), to_signed(1036638064, 32),
     to_signed(1036584389, 32), to_signed(1036530675, 32), to_signed(1036476924, 32), to_signed(1036423135, 32),
     to_signed(1036369307, 32), to_signed(1036315441, 32), to_signed(1036261537, 32), to_signed(1036207595, 32),
     to_signed(1036153615, 32), to_signed(1036099597, 32), to_signed(1036045541, 32), to_signed(1035991447, 32),
     to_signed(1035937314, 32), to_signed(1035883144, 32), to_signed(1035828935, 32), to_signed(1035774689, 32),
     to_signed(1035720404, 32), to_signed(1035666081, 32), to_signed(1035611720, 32), to_signed(1035557321, 32),
     to_signed(1035502884, 32), to_signed(1035448409, 32), to_signed(1035393896, 32), to_signed(1035339345, 32),
     to_signed(1035284755, 32), to_signed(1035230128, 32), to_signed(1035175463, 32), to_signed(1035120759, 32),
     to_signed(1035066018, 32), to_signed(1035011238, 32), to_signed(1034956420, 32), to_signed(1034901565, 32),
     to_signed(1034846671, 32), to_signed(1034791739, 32), to_signed(1034736769, 32), to_signed(1034681761, 32),
     to_signed(1034626715, 32), to_signed(1034571631, 32), to_signed(1034516509, 32), to_signed(1034461349, 32),
     to_signed(1034406151, 32), to_signed(1034350915, 32), to_signed(1034295641, 32), to_signed(1034240329, 32),
     to_signed(1034184978, 32), to_signed(1034129590, 32), to_signed(1034074164, 32), to_signed(1034018700, 32),
     to_signed(1033963197, 32), to_signed(1033907657, 32), to_signed(1033852079, 32), to_signed(1033796462, 32),
     to_signed(1033740808, 32), to_signed(1033685115, 32), to_signed(1033629385, 32), to_signed(1033573617, 32),
     to_signed(1033517810, 32), to_signed(1033461966, 32), to_signed(1033406084, 32), to_signed(1033350163, 32),
     to_signed(1033294205, 32), to_signed(1033238209, 32), to_signed(1033182174, 32), to_signed(1033126102, 32),
     to_signed(1033069992, 32), to_signed(1033013843, 32), to_signed(1032957657, 32), to_signed(1032901433, 32),
     to_signed(1032845170, 32), to_signed(1032788870, 32), to_signed(1032732532, 32), to_signed(1032676156, 32),
     to_signed(1032619742, 32), to_signed(1032563290, 32), to_signed(1032506800, 32), to_signed(1032450272, 32),
     to_signed(1032393706, 32), to_signed(1032337102, 32), to_signed(1032280460, 32), to_signed(1032223780, 32),
     to_signed(1032167062, 32), to_signed(1032110306, 32), to_signed(1032053513, 32), to_signed(1031996681, 32),
     to_signed(1031939812, 32), to_signed(1031882904, 32), to_signed(1031825959, 32), to_signed(1031768975, 32),
     to_signed(1031711954, 32), to_signed(1031654895, 32), to_signed(1031597797, 32), to_signed(1031540662, 32),
     to_signed(1031483489, 32), to_signed(1031426278, 32), to_signed(1031369029, 32), to_signed(1031311742, 32),
     to_signed(1031254418, 32), to_signed(1031197055, 32), to_signed(1031139655, 32), to_signed(1031082216, 32),
     to_signed(1031024740, 32), to_signed(1030967225, 32), to_signed(1030909673, 32), to_signed(1030852083, 32),
     to_signed(1030794455, 32), to_signed(1030736789, 32), to_signed(1030679085, 32), to_signed(1030621344, 32),
     to_signed(1030563564, 32), to_signed(1030505747, 32), to_signed(1030447891, 32), to_signed(1030389998, 32),
     to_signed(1030332067, 32), to_signed(1030274098, 32), to_signed(1030216091, 32), to_signed(1030158046, 32),
     to_signed(1030099963, 32), to_signed(1030041843, 32), to_signed(1029983684, 32), to_signed(1029925488, 32),
     to_signed(1029867254, 32), to_signed(1029808982, 32), to_signed(1029750672, 32), to_signed(1029692324, 32),
     to_signed(1029633939, 32), to_signed(1029575515, 32), to_signed(1029517054, 32), to_signed(1029458555, 32),
     to_signed(1029400018, 32), to_signed(1029341443, 32), to_signed(1029282830, 32), to_signed(1029224180, 32),
     to_signed(1029165491, 32), to_signed(1029106765, 32), to_signed(1029048001, 32), to_signed(1028989199, 32),
     to_signed(1028930359, 32), to_signed(1028871482, 32), to_signed(1028812566, 32), to_signed(1028753613, 32),
     to_signed(1028694622, 32), to_signed(1028635593, 32), to_signed(1028576527, 32), to_signed(1028517422, 32),
     to_signed(1028458280, 32), to_signed(1028399100, 32), to_signed(1028339882, 32), to_signed(1028280626, 32),
     to_signed(1028221332, 32), to_signed(1028162001, 32), to_signed(1028102632, 32), to_signed(1028043225, 32),
     to_signed(1027983780, 32), to_signed(1027924298, 32), to_signed(1027864777, 32), to_signed(1027805219, 32),
     to_signed(1027745623, 32), to_signed(1027685989, 32), to_signed(1027626318, 32), to_signed(1027566609, 32),
     to_signed(1027506862, 32), to_signed(1027447077, 32), to_signed(1027387254, 32), to_signed(1027327394, 32),
     to_signed(1027267495, 32), to_signed(1027207560, 32), to_signed(1027147586, 32), to_signed(1027087574, 32),
     to_signed(1027027525, 32), to_signed(1026967438, 32), to_signed(1026907313, 32), to_signed(1026847151, 32),
     to_signed(1026786951, 32), to_signed(1026726713, 32), to_signed(1026666437, 32), to_signed(1026606123, 32),
     to_signed(1026545772, 32), to_signed(1026485383, 32), to_signed(1026424956, 32), to_signed(1026364492, 32),
     to_signed(1026303990, 32), to_signed(1026243450, 32), to_signed(1026182872, 32), to_signed(1026122256, 32),
     to_signed(1026061603, 32), to_signed(1026000912, 32), to_signed(1025940184, 32), to_signed(1025879418, 32),
     to_signed(1025818614, 32), to_signed(1025757772, 32), to_signed(1025696892, 32), to_signed(1025635975, 32),
     to_signed(1025575020, 32), to_signed(1025514028, 32), to_signed(1025452997, 32), to_signed(1025391929, 32),
     to_signed(1025330824, 32), to_signed(1025269680, 32), to_signed(1025208499, 32), to_signed(1025147280, 32),
     to_signed(1025086024, 32), to_signed(1025024730, 32), to_signed(1024963398, 32), to_signed(1024902028, 32),
     to_signed(1024840621, 32), to_signed(1024779176, 32), to_signed(1024717694, 32), to_signed(1024656173, 32),
     to_signed(1024594615, 32), to_signed(1024533020, 32), to_signed(1024471386, 32), to_signed(1024409716, 32),
     to_signed(1024348007, 32), to_signed(1024286261, 32), to_signed(1024224477, 32), to_signed(1024162655, 32),
     to_signed(1024100796, 32), to_signed(1024038899, 32), to_signed(1023976964, 32), to_signed(1023914992, 32),
     to_signed(1023852982, 32), to_signed(1023790935, 32), to_signed(1023728850, 32), to_signed(1023666727, 32),
     to_signed(1023604567, 32), to_signed(1023542369, 32), to_signed(1023480133, 32), to_signed(1023417860, 32),
     to_signed(1023355549, 32), to_signed(1023293200, 32), to_signed(1023230814, 32), to_signed(1023168390, 32),
     to_signed(1023105929, 32), to_signed(1023043430, 32), to_signed(1022980893, 32), to_signed(1022918319, 32),
     to_signed(1022855707, 32), to_signed(1022793057, 32), to_signed(1022730370, 32), to_signed(1022667646, 32),
     to_signed(1022604883, 32), to_signed(1022542083, 32), to_signed(1022479246, 32), to_signed(1022416371, 32),
     to_signed(1022353458, 32), to_signed(1022290508, 32), to_signed(1022227520, 32), to_signed(1022164495, 32),
     to_signed(1022101432, 32), to_signed(1022038331, 32), to_signed(1021975193, 32), to_signed(1021912017, 32),
     to_signed(1021848804, 32), to_signed(1021785553, 32), to_signed(1021722264, 32), to_signed(1021658938, 32),
     to_signed(1021595575, 32), to_signed(1021532174, 32), to_signed(1021468735, 32), to_signed(1021405259, 32),
     to_signed(1021341745, 32), to_signed(1021278194, 32), to_signed(1021214605, 32), to_signed(1021150978, 32),
     to_signed(1021087314, 32), to_signed(1021023613, 32), to_signed(1020959873, 32), to_signed(1020896097, 32),
     to_signed(1020832283, 32), to_signed(1020768431, 32), to_signed(1020704542, 32), to_signed(1020640615, 32),
     to_signed(1020576651, 32), to_signed(1020512649, 32), to_signed(1020448610, 32), to_signed(1020384533, 32),
     to_signed(1020320418, 32), to_signed(1020256267, 32), to_signed(1020192077, 32), to_signed(1020127850, 32),
     to_signed(1020063586, 32), to_signed(1019999284, 32), to_signed(1019934944, 32), to_signed(1019870568, 32),
     to_signed(1019806153, 32), to_signed(1019741701, 32), to_signed(1019677212, 32), to_signed(1019612685, 32),
     to_signed(1019548121, 32), to_signed(1019483519, 32), to_signed(1019418879, 32), to_signed(1019354203, 32),
     to_signed(1019289488, 32), to_signed(1019224736, 32), to_signed(1019159947, 32), to_signed(1019095120, 32),
     to_signed(1019030256, 32), to_signed(1018965355, 32), to_signed(1018900415, 32), to_signed(1018835439, 32),
     to_signed(1018770425, 32), to_signed(1018705373, 32), to_signed(1018640284, 32), to_signed(1018575158, 32),
     to_signed(1018509994, 32), to_signed(1018444793, 32), to_signed(1018379554, 32), to_signed(1018314278, 32),
     to_signed(1018248964, 32), to_signed(1018183613, 32), to_signed(1018118225, 32), to_signed(1018052799, 32),
     to_signed(1017987335, 32), to_signed(1017921834, 32), to_signed(1017856296, 32), to_signed(1017790720, 32),
     to_signed(1017725107, 32), to_signed(1017659457, 32), to_signed(1017593769, 32), to_signed(1017528044, 32),
     to_signed(1017462281, 32), to_signed(1017396481, 32), to_signed(1017330643, 32), to_signed(1017264768, 32),
     to_signed(1017198856, 32), to_signed(1017132906, 32), to_signed(1017066919, 32), to_signed(1017000894, 32),
     to_signed(1016934832, 32), to_signed(1016868733, 32), to_signed(1016802596, 32), to_signed(1016736422, 32),
     to_signed(1016670211, 32), to_signed(1016603962, 32), to_signed(1016537676, 32), to_signed(1016471352, 32),
     to_signed(1016404991, 32), to_signed(1016338593, 32), to_signed(1016272157, 32), to_signed(1016205684, 32),
     to_signed(1016139173, 32), to_signed(1016072626, 32), to_signed(1016006040, 32), to_signed(1015939418, 32),
     to_signed(1015872758, 32), to_signed(1015806061, 32), to_signed(1015739326, 32), to_signed(1015672554, 32),
     to_signed(1015605745, 32), to_signed(1015538898, 32), to_signed(1015472014, 32), to_signed(1015405093, 32),
     to_signed(1015338134, 32), to_signed(1015271138, 32), to_signed(1015204105, 32), to_signed(1015137034, 32),
     to_signed(1015069927, 32), to_signed(1015002781, 32), to_signed(1014935599, 32), to_signed(1014868379, 32),
     to_signed(1014801122, 32), to_signed(1014733827, 32), to_signed(1014666495, 32), to_signed(1014599126, 32),
     to_signed(1014531720, 32), to_signed(1014464276, 32), to_signed(1014396795, 32), to_signed(1014329277, 32),
     to_signed(1014261721, 32), to_signed(1014194128, 32), to_signed(1014126498, 32), to_signed(1014058830, 32),
     to_signed(1013991126, 32), to_signed(1013923383, 32), to_signed(1013855604, 32), to_signed(1013787787, 32),
     to_signed(1013719934, 32), to_signed(1013652042, 32), to_signed(1013584114, 32), to_signed(1013516148, 32),
     to_signed(1013448145, 32), to_signed(1013380105, 32), to_signed(1013312028, 32), to_signed(1013243913, 32),
     to_signed(1013175761, 32), to_signed(1013107572, 32), to_signed(1013039345, 32), to_signed(1012971081, 32),
     to_signed(1012902780, 32), to_signed(1012834442, 32), to_signed(1012766067, 32), to_signed(1012697654, 32),
     to_signed(1012629204, 32), to_signed(1012560717, 32), to_signed(1012492193, 32), to_signed(1012423631, 32),
     to_signed(1012355032, 32), to_signed(1012286396, 32), to_signed(1012217723, 32), to_signed(1012149012, 32),
     to_signed(1012080264, 32), to_signed(1012011480, 32), to_signed(1011942657, 32), to_signed(1011873798, 32),
     to_signed(1011804901, 32), to_signed(1011735968, 32), to_signed(1011666997, 32), to_signed(1011597989, 32),
     to_signed(1011528943, 32), to_signed(1011459861, 32), to_signed(1011390741, 32), to_signed(1011321584, 32),
     to_signed(1011252390, 32), to_signed(1011183159, 32), to_signed(1011113890, 32), to_signed(1011044585, 32),
     to_signed(1010975242, 32), to_signed(1010905862, 32), to_signed(1010836445, 32), to_signed(1010766991, 32),
     to_signed(1010697499, 32), to_signed(1010627970, 32), to_signed(1010558405, 32), to_signed(1010488802, 32),
     to_signed(1010419162, 32), to_signed(1010349484, 32), to_signed(1010279770, 32), to_signed(1010210018, 32),
     to_signed(1010140230, 32), to_signed(1010070404, 32), to_signed(1010000541, 32), to_signed(1009930641, 32),
     to_signed(1009860704, 32), to_signed(1009790729, 32), to_signed(1009720718, 32), to_signed(1009650669, 32),
     to_signed(1009580584, 32), to_signed(1009510461, 32), to_signed(1009440301, 32), to_signed(1009370104, 32),
     to_signed(1009299870, 32), to_signed(1009229598, 32), to_signed(1009159290, 32), to_signed(1009088944, 32),
     to_signed(1009018562, 32), to_signed(1008948142, 32), to_signed(1008877685, 32), to_signed(1008807191, 32),
     to_signed(1008736660, 32), to_signed(1008666092, 32), to_signed(1008595487, 32), to_signed(1008524845, 32),
     to_signed(1008454166, 32), to_signed(1008383449, 32), to_signed(1008312696, 32), to_signed(1008241905, 32),
     to_signed(1008171077, 32), to_signed(1008100213, 32), to_signed(1008029311, 32), to_signed(1007958372, 32),
     to_signed(1007887396, 32), to_signed(1007816383, 32), to_signed(1007745333, 32), to_signed(1007674246, 32),
     to_signed(1007603122, 32), to_signed(1007531961, 32), to_signed(1007460763, 32), to_signed(1007389528, 32),
     to_signed(1007318256, 32), to_signed(1007246946, 32), to_signed(1007175600, 32), to_signed(1007104217, 32),
     to_signed(1007032796, 32), to_signed(1006961339, 32), to_signed(1006889844, 32), to_signed(1006818313, 32),
     to_signed(1006746744, 32), to_signed(1006675139, 32), to_signed(1006603496, 32), to_signed(1006531817, 32),
     to_signed(1006460100, 32), to_signed(1006388347, 32), to_signed(1006316556, 32), to_signed(1006244729, 32),
     to_signed(1006172864, 32), to_signed(1006100963, 32), to_signed(1006029024, 32), to_signed(1005957049, 32),
     to_signed(1005885036, 32), to_signed(1005812987, 32), to_signed(1005740900, 32), to_signed(1005668777, 32),
     to_signed(1005596617, 32), to_signed(1005524419, 32), to_signed(1005452185, 32), to_signed(1005379913, 32),
     to_signed(1005307605, 32), to_signed(1005235260, 32), to_signed(1005162878, 32), to_signed(1005090459, 32),
     to_signed(1005018003, 32), to_signed(1004945509, 32), to_signed(1004872979, 32), to_signed(1004800412, 32),
     to_signed(1004727809, 32), to_signed(1004655168, 32), to_signed(1004582490, 32), to_signed(1004509775, 32),
     to_signed(1004437024, 32), to_signed(1004364235, 32), to_signed(1004291410, 32), to_signed(1004218547, 32),
     to_signed(1004145648, 32), to_signed(1004072711, 32), to_signed(1003999738, 32), to_signed(1003926728, 32),
     to_signed(1003853681, 32), to_signed(1003780597, 32), to_signed(1003707476, 32), to_signed(1003634319, 32),
     to_signed(1003561124, 32), to_signed(1003487893, 32), to_signed(1003414624, 32), to_signed(1003341319, 32),
     to_signed(1003267977, 32), to_signed(1003194597, 32), to_signed(1003121181, 32), to_signed(1003047729, 32),
     to_signed(1002974239, 32), to_signed(1002900712, 32), to_signed(1002827149, 32), to_signed(1002753548, 32),
     to_signed(1002679911, 32), to_signed(1002606237, 32), to_signed(1002532526, 32), to_signed(1002458778, 32),
     to_signed(1002384994, 32), to_signed(1002311172, 32), to_signed(1002237314, 32), to_signed(1002163418, 32),
     to_signed(1002089486, 32), to_signed(1002015517, 32), to_signed(1001941512, 32), to_signed(1001867469, 32),
     to_signed(1001793390, 32), to_signed(1001719273, 32), to_signed(1001645120, 32), to_signed(1001570930, 32),
     to_signed(1001496704, 32), to_signed(1001422440, 32), to_signed(1001348140, 32), to_signed(1001273802, 32),
     to_signed(1001199428, 32), to_signed(1001125017, 32), to_signed(1001050570, 32), to_signed(1000976085, 32),
     to_signed(1000901564, 32), to_signed(1000827006, 32), to_signed(1000752411, 32), to_signed(1000677780, 32),
     to_signed(1000603111, 32), to_signed(1000528406, 32), to_signed(1000453664, 32), to_signed(1000378885, 32),
     to_signed(1000304069, 32), to_signed(1000229217, 32), to_signed(1000154328, 32), to_signed(1000079402, 32),
     to_signed(1000004439, 32), to_signed(999929440, 32), to_signed(999854404, 32), to_signed(999779331, 32),
     to_signed(999704221, 32), to_signed(999629074, 32), to_signed(999553891, 32), to_signed(999478671, 32),
     to_signed(999403415, 32), to_signed(999328121, 32), to_signed(999252791, 32), to_signed(999177424, 32),
     to_signed(999102020, 32), to_signed(999026580, 32), to_signed(998951103, 32), to_signed(998875589, 32),
     to_signed(998800038, 32), to_signed(998724451, 32), to_signed(998648827, 32), to_signed(998573166, 32),
     to_signed(998497468, 32), to_signed(998421734, 32), to_signed(998345963, 32), to_signed(998270156, 32),
     to_signed(998194311, 32), to_signed(998118430, 32), to_signed(998042512, 32), to_signed(997966558, 32),
     to_signed(997890567, 32), to_signed(997814539, 32), to_signed(997738475, 32), to_signed(997662373, 32),
     to_signed(997586236, 32), to_signed(997510061, 32), to_signed(997433850, 32), to_signed(997357602, 32),
     to_signed(997281317, 32), to_signed(997204996, 32), to_signed(997128638, 32), to_signed(997052244, 32),
     to_signed(996975812, 32), to_signed(996899345, 32), to_signed(996822840, 32), to_signed(996746299, 32),
     to_signed(996669721, 32), to_signed(996593107, 32), to_signed(996516456, 32), to_signed(996439768, 32),
     to_signed(996363043, 32), to_signed(996286282, 32), to_signed(996209485, 32), to_signed(996132650, 32),
     to_signed(996055780, 32), to_signed(995978872, 32), to_signed(995901928, 32), to_signed(995824947, 32),
     to_signed(995747930, 32), to_signed(995670876, 32), to_signed(995593785, 32), to_signed(995516658, 32),
     to_signed(995439494, 32), to_signed(995362294, 32), to_signed(995285057, 32), to_signed(995207783, 32),
     to_signed(995130473, 32), to_signed(995053126, 32), to_signed(994975743, 32), to_signed(994898323, 32),
     to_signed(994820867, 32), to_signed(994743373, 32), to_signed(994665844, 32), to_signed(994588278, 32),
     to_signed(994510675, 32), to_signed(994433035, 32), to_signed(994355360, 32), to_signed(994277647, 32),
     to_signed(994199898, 32), to_signed(994122112, 32), to_signed(994044290, 32), to_signed(993966432, 32),
     to_signed(993888536, 32), to_signed(993810605, 32), to_signed(993732636, 32), to_signed(993654631, 32),
     to_signed(993576590, 32), to_signed(993498512, 32), to_signed(993420398, 32), to_signed(993342247, 32),
     to_signed(993264059, 32), to_signed(993185835, 32), to_signed(993107575, 32), to_signed(993029277, 32),
     to_signed(992950944, 32), to_signed(992872574, 32), to_signed(992794167, 32), to_signed(992715724, 32),
     to_signed(992637245, 32), to_signed(992558729, 32), to_signed(992480176, 32), to_signed(992401587, 32),
     to_signed(992322961, 32), to_signed(992244299, 32), to_signed(992165601, 32), to_signed(992086866, 32),
     to_signed(992008094, 32), to_signed(991929286, 32), to_signed(991850442, 32), to_signed(991771561, 32),
     to_signed(991692644, 32), to_signed(991613690, 32), to_signed(991534700, 32), to_signed(991455673, 32),
     to_signed(991376610, 32), to_signed(991297510, 32), to_signed(991218374, 32), to_signed(991139202, 32),
     to_signed(991059993, 32), to_signed(990980747, 32), to_signed(990901465, 32), to_signed(990822147, 32),
     to_signed(990742793, 32), to_signed(990663401, 32), to_signed(990583974, 32), to_signed(990504510, 32),
     to_signed(990425010, 32), to_signed(990345473, 32), to_signed(990265900, 32), to_signed(990186290, 32),
     to_signed(990106644, 32), to_signed(990026961, 32), to_signed(989947243, 32), to_signed(989867487, 32),
     to_signed(989787696, 32), to_signed(989707868, 32), to_signed(989628003, 32), to_signed(989548103, 32),
     to_signed(989468165, 32), to_signed(989388192, 32), to_signed(989308182, 32), to_signed(989228136, 32),
     to_signed(989148053, 32), to_signed(989067934, 32), to_signed(988987779, 32), to_signed(988907587, 32),
     to_signed(988827359, 32), to_signed(988747094, 32), to_signed(988666793, 32), to_signed(988586456, 32),
     to_signed(988506083, 32), to_signed(988425673, 32), to_signed(988345227, 32), to_signed(988264744, 32),
     to_signed(988184225, 32), to_signed(988103670, 32), to_signed(988023078, 32), to_signed(987942450, 32),
     to_signed(987861786, 32), to_signed(987781086, 32), to_signed(987700349, 32), to_signed(987619576, 32),
     to_signed(987538766, 32), to_signed(987457920, 32), to_signed(987377038, 32), to_signed(987296120, 32),
     to_signed(987215165, 32), to_signed(987134174, 32), to_signed(987053147, 32), to_signed(986972083, 32),
     to_signed(986890984, 32), to_signed(986809847, 32), to_signed(986728675, 32), to_signed(986647466, 32),
     to_signed(986566221, 32), to_signed(986484940, 32), to_signed(986403623, 32), to_signed(986322269, 32),
     to_signed(986240879, 32), to_signed(986159452, 32), to_signed(986077990, 32), to_signed(985996491, 32),
     to_signed(985914956, 32), to_signed(985833385, 32), to_signed(985751777, 32), to_signed(985670133, 32),
     to_signed(985588453, 32), to_signed(985506737, 32), to_signed(985424984, 32), to_signed(985343195, 32),
     to_signed(985261370, 32), to_signed(985179509, 32), to_signed(985097612, 32), to_signed(985015678, 32),
     to_signed(984933708, 32), to_signed(984851702, 32), to_signed(984769660, 32), to_signed(984687581, 32),
     to_signed(984605467, 32), to_signed(984523316, 32), to_signed(984441129, 32), to_signed(984358905, 32),
     to_signed(984276646, 32), to_signed(984194350, 32), to_signed(984112018, 32), to_signed(984029650, 32),
     to_signed(983947246, 32), to_signed(983864806, 32), to_signed(983782329, 32), to_signed(983699816, 32),
     to_signed(983617267, 32), to_signed(983534682, 32), to_signed(983452061, 32), to_signed(983369404, 32),
     to_signed(983286710, 32), to_signed(983203980, 32), to_signed(983121214, 32), to_signed(983038412, 32),
     to_signed(982955574, 32), to_signed(982872700, 32), to_signed(982789789, 32), to_signed(982706843, 32),
     to_signed(982623860, 32), to_signed(982540841, 32), to_signed(982457786, 32), to_signed(982374695, 32),
     to_signed(982291568, 32), to_signed(982208405, 32), to_signed(982125205, 32), to_signed(982041970, 32),
     to_signed(981958698, 32), to_signed(981875390, 32), to_signed(981792047, 32), to_signed(981708667, 32),
     to_signed(981625251, 32), to_signed(981541798, 32), to_signed(981458310, 32), to_signed(981374786, 32),
     to_signed(981291226, 32), to_signed(981207629, 32), to_signed(981123997, 32), to_signed(981040328, 32),
     to_signed(980956623, 32), to_signed(980872882, 32), to_signed(980789106, 32), to_signed(980705293, 32),
     to_signed(980621444, 32), to_signed(980537559, 32), to_signed(980453638, 32), to_signed(980369681, 32),
     to_signed(980285688, 32), to_signed(980201658, 32), to_signed(980117593, 32), to_signed(980033492, 32),
     to_signed(979949355, 32), to_signed(979865181, 32), to_signed(979780972, 32), to_signed(979696727, 32),
     to_signed(979612445, 32), to_signed(979528128, 32), to_signed(979443774, 32), to_signed(979359385, 32),
     to_signed(979274960, 32), to_signed(979190498, 32), to_signed(979106001, 32), to_signed(979021467, 32),
     to_signed(978936898, 32), to_signed(978852292, 32), to_signed(978767651, 32), to_signed(978682973, 32),
     to_signed(978598260, 32), to_signed(978513511, 32), to_signed(978428725, 32), to_signed(978343904, 32),
     to_signed(978259047, 32), to_signed(978174153, 32), to_signed(978089224, 32), to_signed(978004259, 32),
     to_signed(977919258, 32), to_signed(977834221, 32), to_signed(977749148, 32), to_signed(977664039, 32),
     to_signed(977578894, 32), to_signed(977493713, 32), to_signed(977408496, 32), to_signed(977323243, 32),
     to_signed(977237955, 32), to_signed(977152630, 32), to_signed(977067269, 32), to_signed(976981873, 32),
     to_signed(976896441, 32), to_signed(976810972, 32), to_signed(976725468, 32), to_signed(976639928, 32),
     to_signed(976554352, 32), to_signed(976468740, 32), to_signed(976383092, 32), to_signed(976297408, 32),
     to_signed(976211688, 32), to_signed(976125933, 32), to_signed(976040141, 32), to_signed(975954314, 32),
     to_signed(975868451, 32), to_signed(975782552, 32), to_signed(975696617, 32), to_signed(975610646, 32),
     to_signed(975524639, 32), to_signed(975438597, 32), to_signed(975352518, 32), to_signed(975266404, 32),
     to_signed(975180254, 32), to_signed(975094068, 32), to_signed(975007846, 32), to_signed(974921588, 32),
     to_signed(974835295, 32), to_signed(974748965, 32), to_signed(974662600, 32), to_signed(974576199, 32),
     to_signed(974489762, 32), to_signed(974403289, 32), to_signed(974316781, 32), to_signed(974230236, 32),
     to_signed(974143656, 32), to_signed(974057040, 32), to_signed(973970388, 32), to_signed(973883701, 32),
     to_signed(973796977, 32), to_signed(973710218, 32), to_signed(973623423, 32), to_signed(973536592, 32),
     to_signed(973449725, 32), to_signed(973362823, 32), to_signed(973275885, 32), to_signed(973188911, 32),
     to_signed(973101901, 32), to_signed(973014855, 32), to_signed(972927774, 32), to_signed(972840657, 32),
     to_signed(972753504, 32), to_signed(972666315, 32), to_signed(972579091, 32), to_signed(972491831, 32),
     to_signed(972404535, 32), to_signed(972317203, 32), to_signed(972229836, 32), to_signed(972142433, 32),
     to_signed(972054994, 32), to_signed(971967519, 32), to_signed(971880009, 32), to_signed(971792462, 32),
     to_signed(971704881, 32), to_signed(971617263, 32), to_signed(971529610, 32), to_signed(971441921, 32),
     to_signed(971354196, 32), to_signed(971266435, 32), to_signed(971178639, 32), to_signed(971090807, 32),
     to_signed(971002940, 32), to_signed(970915037, 32), to_signed(970827098, 32), to_signed(970739123, 32),
     to_signed(970651112, 32), to_signed(970563066, 32), to_signed(970474985, 32), to_signed(970386867, 32),
     to_signed(970298714, 32), to_signed(970210525, 32), to_signed(970122301, 32), to_signed(970034041, 32),
     to_signed(969945745, 32), to_signed(969857414, 32), to_signed(969769046, 32), to_signed(969680644, 32),
     to_signed(969592205, 32), to_signed(969503731, 32), to_signed(969415222, 32), to_signed(969326676, 32),
     to_signed(969238095, 32), to_signed(969149479, 32), to_signed(969060826, 32), to_signed(968972138, 32),
     to_signed(968883415, 32), to_signed(968794656, 32), to_signed(968705861, 32), to_signed(968617031, 32),
     to_signed(968528165, 32), to_signed(968439263, 32), to_signed(968350326, 32), to_signed(968261353, 32),
     to_signed(968172345, 32), to_signed(968083301, 32), to_signed(967994221, 32), to_signed(967905106, 32),
     to_signed(967815955, 32), to_signed(967726769, 32), to_signed(967637547, 32), to_signed(967548289, 32),
     to_signed(967458996, 32), to_signed(967369668, 32), to_signed(967280303, 32), to_signed(967190904, 32),
     to_signed(967101468, 32), to_signed(967011997, 32), to_signed(966922491, 32), to_signed(966832949, 32),
     to_signed(966743371, 32), to_signed(966653758, 32), to_signed(966564109, 32), to_signed(966474425, 32),
     to_signed(966384706, 32), to_signed(966294950, 32), to_signed(966205159, 32), to_signed(966115333, 32),
     to_signed(966025471, 32), to_signed(965935574, 32), to_signed(965845641, 32), to_signed(965755673, 32),
     to_signed(965665669, 32), to_signed(965575630, 32), to_signed(965485555, 32), to_signed(965395444, 32),
     to_signed(965305298, 32), to_signed(965215117, 32), to_signed(965124900, 32), to_signed(965034648, 32),
     to_signed(964944360, 32), to_signed(964854037, 32), to_signed(964763678, 32), to_signed(964673284, 32),
     to_signed(964582854, 32), to_signed(964492389, 32), to_signed(964401888, 32), to_signed(964311352, 32),
     to_signed(964220780, 32), to_signed(964130173, 32), to_signed(964039531, 32), to_signed(963948853, 32),
     to_signed(963858140, 32), to_signed(963767391, 32), to_signed(963676607, 32), to_signed(963585787, 32),
     to_signed(963494932, 32), to_signed(963404042, 32), to_signed(963313116, 32), to_signed(963222154, 32),
     to_signed(963131157, 32), to_signed(963040125, 32), to_signed(962949058, 32), to_signed(962857955, 32),
     to_signed(962766816, 32), to_signed(962675643, 32), to_signed(962584433, 32), to_signed(962493189, 32),
     to_signed(962401909, 32), to_signed(962310594, 32), to_signed(962219243, 32), to_signed(962127857, 32),
     to_signed(962036435, 32), to_signed(961944978, 32), to_signed(961853486, 32), to_signed(961761959, 32),
     to_signed(961670396, 32), to_signed(961578797, 32), to_signed(961487164, 32), to_signed(961395495, 32),
     to_signed(961303790, 32), to_signed(961212051, 32), to_signed(961120276, 32), to_signed(961028465, 32),
     to_signed(960936620, 32), to_signed(960844739, 32), to_signed(960752822, 32), to_signed(960660870, 32),
     to_signed(960568883, 32), to_signed(960476861, 32), to_signed(960384803, 32), to_signed(960292711, 32),
     to_signed(960200582, 32), to_signed(960108419, 32), to_signed(960016220, 32), to_signed(959923986, 32),
     to_signed(959831716, 32), to_signed(959739411, 32), to_signed(959647071, 32), to_signed(959554696, 32),
     to_signed(959462286, 32), to_signed(959369840, 32), to_signed(959277359, 32), to_signed(959184842, 32),
     to_signed(959092290, 32), to_signed(958999703, 32), to_signed(958907081, 32), to_signed(958814424, 32),
     to_signed(958721731, 32), to_signed(958629003, 32), to_signed(958536240, 32), to_signed(958443441, 32),
     to_signed(958350608, 32), to_signed(958257739, 32), to_signed(958164835, 32), to_signed(958071895, 32),
     to_signed(957978921, 32), to_signed(957885911, 32), to_signed(957792866, 32), to_signed(957699786, 32),
     to_signed(957606670, 32), to_signed(957513519, 32), to_signed(957420333, 32), to_signed(957327112, 32),
     to_signed(957233856, 32), to_signed(957140565, 32), to_signed(957047238, 32), to_signed(956953876, 32),
     to_signed(956860479, 32), to_signed(956767047, 32), to_signed(956673579, 32), to_signed(956580077, 32),
     to_signed(956486539, 32), to_signed(956392966, 32), to_signed(956299358, 32), to_signed(956205715, 32),
     to_signed(956112036, 32), to_signed(956018323, 32), to_signed(955924574, 32), to_signed(955830790, 32),
     to_signed(955736971, 32), to_signed(955643117, 32), to_signed(955549228, 32), to_signed(955455303, 32),
     to_signed(955361344, 32), to_signed(955267349, 32), to_signed(955173319, 32), to_signed(955079254, 32),
     to_signed(954985154, 32), to_signed(954891019, 32), to_signed(954796849, 32), to_signed(954702644, 32),
     to_signed(954608403, 32), to_signed(954514128, 32), to_signed(954419817, 32), to_signed(954325471, 32),
     to_signed(954231090, 32), to_signed(954136675, 32), to_signed(954042224, 32), to_signed(953947738, 32),
     to_signed(953853216, 32), to_signed(953758660, 32), to_signed(953664069, 32), to_signed(953569443, 32),
     to_signed(953474781, 32), to_signed(953380085, 32), to_signed(953285353, 32), to_signed(953190587, 32),
     to_signed(953095785, 32), to_signed(953000948, 32), to_signed(952906077, 32), to_signed(952811170, 32),
     to_signed(952716228, 32), to_signed(952621251, 32), to_signed(952526240, 32), to_signed(952431193, 32),
     to_signed(952336111, 32), to_signed(952240994, 32), to_signed(952145842, 32), to_signed(952050655, 32),
     to_signed(951955434, 32), to_signed(951860177, 32), to_signed(951764885, 32), to_signed(951669558, 32),
     to_signed(951574196, 32), to_signed(951478799, 32), to_signed(951383367, 32), to_signed(951287900, 32),
     to_signed(951192399, 32), to_signed(951096862, 32), to_signed(951001290, 32), to_signed(950905684, 32),
     to_signed(950810042, 32), to_signed(950714365, 32), to_signed(950618654, 32), to_signed(950522907, 32),
     to_signed(950427126, 32), to_signed(950331309, 32), to_signed(950235458, 32), to_signed(950139572, 32),
     to_signed(950043650, 32), to_signed(949947694, 32), to_signed(949851703, 32), to_signed(949755677, 32),
     to_signed(949659616, 32), to_signed(949563520, 32), to_signed(949467390, 32), to_signed(949371224, 32),
     to_signed(949275023, 32), to_signed(949178788, 32), to_signed(949082517, 32), to_signed(948986212, 32),
     to_signed(948889872, 32), to_signed(948793497, 32), to_signed(948697087, 32), to_signed(948600642, 32),
     to_signed(948504163, 32), to_signed(948407648, 32), to_signed(948311099, 32), to_signed(948214514, 32),
     to_signed(948117895, 32), to_signed(948021241, 32), to_signed(947924552, 32), to_signed(947827828, 32),
     to_signed(947731070, 32), to_signed(947634276, 32), to_signed(947537448, 32), to_signed(947440585, 32),
     to_signed(947343687, 32), to_signed(947246754, 32), to_signed(947149787, 32), to_signed(947052784, 32),
     to_signed(946955747, 32), to_signed(946858675, 32), to_signed(946761568, 32), to_signed(946664426, 32),
     to_signed(946567250, 32), to_signed(946470039, 32), to_signed(946372792, 32), to_signed(946275512, 32),
     to_signed(946178196, 32), to_signed(946080845, 32), to_signed(945983460, 32), to_signed(945886040, 32),
     to_signed(945788585, 32), to_signed(945691096, 32), to_signed(945593571, 32), to_signed(945496012, 32),
     to_signed(945398418, 32), to_signed(945300790, 32), to_signed(945203126, 32), to_signed(945105428, 32),
     to_signed(945007695, 32), to_signed(944909928, 32), to_signed(944812125, 32), to_signed(944714288, 32),
     to_signed(944616416, 32), to_signed(944518510, 32), to_signed(944420568, 32), to_signed(944322592, 32),
     to_signed(944224582, 32), to_signed(944126536, 32), to_signed(944028456, 32), to_signed(943930341, 32),
     to_signed(943832191, 32), to_signed(943734007, 32), to_signed(943635788, 32), to_signed(943537534, 32),
     to_signed(943439246, 32), to_signed(943340923, 32), to_signed(943242565, 32), to_signed(943144173, 32),
     to_signed(943045745, 32), to_signed(942947284, 32), to_signed(942848787, 32), to_signed(942750256, 32),
     to_signed(942651690, 32), to_signed(942553090, 32), to_signed(942454455, 32), to_signed(942355785, 32),
     to_signed(942257081, 32), to_signed(942158341, 32), to_signed(942059568, 32), to_signed(941960759, 32),
     to_signed(941861917, 32), to_signed(941763039, 32), to_signed(941664127, 32), to_signed(941565180, 32),
     to_signed(941466198, 32), to_signed(941367182, 32), to_signed(941268132, 32), to_signed(941169046, 32),
     to_signed(941069926, 32), to_signed(940970772, 32), to_signed(940871583, 32), to_signed(940772359, 32),
     to_signed(940673101, 32), to_signed(940573808, 32), to_signed(940474481, 32), to_signed(940375119, 32),
     to_signed(940275722, 32), to_signed(940176291, 32), to_signed(940076825, 32), to_signed(939977325, 32),
     to_signed(939877790, 32), to_signed(939778220, 32), to_signed(939678616, 32), to_signed(939578978, 32),
     to_signed(939479305, 32), to_signed(939379597, 32), to_signed(939279855, 32), to_signed(939180078, 32),
     to_signed(939080267, 32), to_signed(938980422, 32), to_signed(938880541, 32), to_signed(938780626, 32),
     to_signed(938680677, 32), to_signed(938580693, 32), to_signed(938480675, 32), to_signed(938380622, 32),
     to_signed(938280535, 32), to_signed(938180413, 32), to_signed(938080257, 32), to_signed(937980066, 32),
     to_signed(937879841, 32), to_signed(937779581, 32), to_signed(937679287, 32), to_signed(937578958, 32),
     to_signed(937478595, 32), to_signed(937378197, 32), to_signed(937277765, 32), to_signed(937177298, 32),
     to_signed(937076797, 32), to_signed(936976262, 32), to_signed(936875692, 32), to_signed(936775087, 32),
     to_signed(936674448, 32), to_signed(936573775, 32), to_signed(936473067, 32), to_signed(936372325, 32),
     to_signed(936271549, 32), to_signed(936170738, 32), to_signed(936069892, 32), to_signed(935969012, 32),
     to_signed(935868098, 32), to_signed(935767149, 32), to_signed(935666166, 32), to_signed(935565149, 32),
     to_signed(935464097, 32), to_signed(935363011, 32), to_signed(935261890, 32), to_signed(935160735, 32),
     to_signed(935059546, 32), to_signed(934958322, 32), to_signed(934857064, 32), to_signed(934755771, 32),
     to_signed(934654444, 32), to_signed(934553083, 32), to_signed(934451687, 32), to_signed(934350257, 32),
     to_signed(934248793, 32), to_signed(934147294, 32), to_signed(934045761, 32), to_signed(933944194, 32),
     to_signed(933842592, 32), to_signed(933740956, 32), to_signed(933639286, 32), to_signed(933537581, 32),
     to_signed(933435842, 32), to_signed(933334068, 32), to_signed(933232261, 32), to_signed(933130419, 32),
     to_signed(933028542, 32), to_signed(932926632, 32), to_signed(932824687, 32), to_signed(932722708, 32),
     to_signed(932620694, 32), to_signed(932518646, 32), to_signed(932416564, 32), to_signed(932314448, 32),
     to_signed(932212297, 32), to_signed(932110112, 32), to_signed(932007893, 32), to_signed(931905640, 32),
     to_signed(931803352, 32), to_signed(931701030, 32), to_signed(931598674, 32), to_signed(931496283, 32),
     to_signed(931393859, 32), to_signed(931291400, 32), to_signed(931188906, 32), to_signed(931086379, 32),
     to_signed(930983817, 32), to_signed(930881221, 32), to_signed(930778591, 32), to_signed(930675927, 32),
     to_signed(930573228, 32), to_signed(930470495, 32), to_signed(930367728, 32), to_signed(930264927, 32),
     to_signed(930162092, 32), to_signed(930059222, 32), to_signed(929956318, 32), to_signed(929853380, 32),
     to_signed(929750408, 32), to_signed(929647402, 32), to_signed(929544361, 32), to_signed(929441286, 32),
     to_signed(929338177, 32), to_signed(929235034, 32), to_signed(929131857, 32), to_signed(929028646, 32),
     to_signed(928925400, 32), to_signed(928822120, 32), to_signed(928718807, 32), to_signed(928615459, 32),
     to_signed(928512076, 32), to_signed(928408660, 32), to_signed(928305210, 32), to_signed(928201725, 32),
     to_signed(928098206, 32), to_signed(927994654, 32), to_signed(927891067, 32), to_signed(927787446, 32),
     to_signed(927683790, 32), to_signed(927580101, 32), to_signed(927476378, 32), to_signed(927372620, 32),
     to_signed(927268829, 32), to_signed(927165003, 32), to_signed(927061143, 32), to_signed(926957249, 32),
     to_signed(926853322, 32), to_signed(926749360, 32), to_signed(926645363, 32), to_signed(926541333, 32),
     to_signed(926437269, 32), to_signed(926333171, 32), to_signed(926229039, 32), to_signed(926124872, 32),
     to_signed(926020672, 32), to_signed(925916437, 32), to_signed(925812169, 32), to_signed(925707866, 32),
     to_signed(925603530, 32), to_signed(925499159, 32), to_signed(925394754, 32), to_signed(925290316, 32),
     to_signed(925185843, 32), to_signed(925081336, 32), to_signed(924976795, 32), to_signed(924872221, 32),
     to_signed(924767612, 32), to_signed(924662969, 32), to_signed(924558292, 32), to_signed(924453582, 32),
     to_signed(924348837, 32), to_signed(924244058, 32), to_signed(924139246, 32), to_signed(924034399, 32),
     to_signed(923929518, 32), to_signed(923824604, 32), to_signed(923719655, 32), to_signed(923614672, 32),
     to_signed(923509656, 32), to_signed(923404605, 32), to_signed(923299521, 32), to_signed(923194403, 32),
     to_signed(923089250, 32), to_signed(922984064, 32), to_signed(922878844, 32), to_signed(922773590, 32),
     to_signed(922668302, 32), to_signed(922562980, 32), to_signed(922457624, 32), to_signed(922352234, 32),
     to_signed(922246810, 32), to_signed(922141353, 32), to_signed(922035861, 32), to_signed(921930336, 32),
     to_signed(921824777, 32), to_signed(921719183, 32), to_signed(921613556, 32), to_signed(921507895, 32),
     to_signed(921402200, 32), to_signed(921296472, 32), to_signed(921190709, 32), to_signed(921084913, 32),
     to_signed(920979082, 32), to_signed(920873218, 32), to_signed(920767320, 32), to_signed(920661388, 32),
     to_signed(920555422, 32), to_signed(920449423, 32), to_signed(920343389, 32), to_signed(920237322, 32),
     to_signed(920131221, 32), to_signed(920025086, 32), to_signed(919918917, 32), to_signed(919812714, 32),
     to_signed(919706478, 32), to_signed(919600208, 32), to_signed(919493904, 32), to_signed(919387566, 32),
     to_signed(919281194, 32), to_signed(919174789, 32), to_signed(919068349, 32), to_signed(918961876, 32),
     to_signed(918855369, 32), to_signed(918748829, 32), to_signed(918642254, 32), to_signed(918535646, 32),
     to_signed(918429004, 32), to_signed(918322328, 32), to_signed(918215619, 32), to_signed(918108876, 32),
     to_signed(918002099, 32), to_signed(917895288, 32), to_signed(917788443, 32), to_signed(917681565, 32),
     to_signed(917574653, 32), to_signed(917467707, 32), to_signed(917360728, 32), to_signed(917253715, 32),
     to_signed(917146668, 32), to_signed(917039587, 32), to_signed(916932473, 32), to_signed(916825325, 32),
     to_signed(916718143, 32), to_signed(916610928, 32), to_signed(916503678, 32), to_signed(916396395, 32),
     to_signed(916289079, 32), to_signed(916181729, 32), to_signed(916074345, 32), to_signed(915966927, 32),
     to_signed(915859476, 32), to_signed(915751991, 32), to_signed(915644472, 32), to_signed(915536920, 32),
     to_signed(915429334, 32), to_signed(915321714, 32), to_signed(915214061, 32), to_signed(915106374, 32),
     to_signed(914998653, 32), to_signed(914890899, 32), to_signed(914783111, 32), to_signed(914675290, 32),
     to_signed(914567435, 32), to_signed(914459546, 32), to_signed(914351624, 32), to_signed(914243668, 32),
     to_signed(914135678, 32), to_signed(914027655, 32), to_signed(913919598, 32), to_signed(913811507, 32),
     to_signed(913703383, 32), to_signed(913595226, 32), to_signed(913487035, 32), to_signed(913378810, 32),
     to_signed(913270551, 32), to_signed(913162259, 32), to_signed(913053934, 32), to_signed(912945575, 32),
     to_signed(912837182, 32), to_signed(912728756, 32), to_signed(912620296, 32), to_signed(912511803, 32),
     to_signed(912403276, 32), to_signed(912294715, 32), to_signed(912186121, 32), to_signed(912077494, 32),
     to_signed(911968833, 32), to_signed(911860138, 32), to_signed(911751410, 32), to_signed(911642649, 32),
     to_signed(911533853, 32), to_signed(911425025, 32), to_signed(911316163, 32), to_signed(911207267, 32),
     to_signed(911098338, 32), to_signed(910989375, 32), to_signed(910880379, 32), to_signed(910771349, 32),
     to_signed(910662286, 32), to_signed(910553189, 32), to_signed(910444059, 32), to_signed(910334896, 32),
     to_signed(910225699, 32), to_signed(910116468, 32), to_signed(910007204, 32), to_signed(909897907, 32),
     to_signed(909788576, 32), to_signed(909679211, 32), to_signed(909569814, 32), to_signed(909460382, 32),
     to_signed(909350918, 32), to_signed(909241420, 32), to_signed(909131888, 32), to_signed(909022323, 32),
     to_signed(908912725, 32), to_signed(908803093, 32), to_signed(908693428, 32), to_signed(908583729, 32),
     to_signed(908473997, 32), to_signed(908364231, 32), to_signed(908254433, 32), to_signed(908144600, 32),
     to_signed(908034735, 32), to_signed(907924836, 32), to_signed(907814903, 32), to_signed(907704938, 32),
     to_signed(907594938, 32), to_signed(907484906, 32), to_signed(907374840, 32), to_signed(907264741, 32),
     to_signed(907154608, 32), to_signed(907044442, 32), to_signed(906934243, 32), to_signed(906824010, 32),
     to_signed(906713744, 32), to_signed(906603445, 32), to_signed(906493112, 32), to_signed(906382746, 32),
     to_signed(906272347, 32), to_signed(906161914, 32), to_signed(906051448, 32), to_signed(905940949, 32),
     to_signed(905830417, 32), to_signed(905719851, 32), to_signed(905609251, 32), to_signed(905498619, 32),
     to_signed(905387953, 32), to_signed(905277254, 32), to_signed(905166522, 32), to_signed(905055756, 32),
     to_signed(904944957, 32), to_signed(904834125, 32), to_signed(904723260, 32), to_signed(904612361, 32),
     to_signed(904501429, 32), to_signed(904390464, 32), to_signed(904279465, 32), to_signed(904168434, 32),
     to_signed(904057369, 32), to_signed(903946270, 32), to_signed(903835139, 32), to_signed(903723974, 32),
     to_signed(903612776, 32), to_signed(903501545, 32), to_signed(903390281, 32), to_signed(903278983, 32),
     to_signed(903167653, 32), to_signed(903056289, 32), to_signed(902944892, 32), to_signed(902833461, 32),
     to_signed(902721998, 32), to_signed(902610501, 32), to_signed(902498971, 32), to_signed(902387408, 32),
     to_signed(902275811, 32), to_signed(902164182, 32), to_signed(902052519, 32), to_signed(901940824, 32),
     to_signed(901829095, 32), to_signed(901717332, 32), to_signed(901605537, 32), to_signed(901493709, 32),
     to_signed(901381847, 32), to_signed(901269952, 32), to_signed(901158025, 32), to_signed(901046064, 32),
     to_signed(900934069, 32), to_signed(900822042, 32), to_signed(900709982, 32), to_signed(900597888, 32),
     to_signed(900485762, 32), to_signed(900373602, 32), to_signed(900261409, 32), to_signed(900149183, 32),
     to_signed(900036924, 32), to_signed(899924632, 32), to_signed(899812307, 32), to_signed(899699949, 32),
     to_signed(899587557, 32), to_signed(899475133, 32), to_signed(899362675, 32), to_signed(899250185, 32),
     to_signed(899137661, 32), to_signed(899025105, 32), to_signed(898912515, 32), to_signed(898799892, 32),
     to_signed(898687236, 32), to_signed(898574547, 32), to_signed(898461825, 32), to_signed(898349070, 32),
     to_signed(898236282, 32), to_signed(898123461, 32), to_signed(898010607, 32), to_signed(897897720, 32),
     to_signed(897784800, 32), to_signed(897671847, 32), to_signed(897558861, 32), to_signed(897445842, 32),
     to_signed(897332790, 32), to_signed(897219705, 32), to_signed(897106587, 32), to_signed(896993436, 32),
     to_signed(896880252, 32), to_signed(896767035, 32), to_signed(896653785, 32), to_signed(896540502, 32),
     to_signed(896427186, 32), to_signed(896313837, 32), to_signed(896200456, 32), to_signed(896087041, 32),
     to_signed(895973593, 32), to_signed(895860112, 32), to_signed(895746599, 32), to_signed(895633052, 32),
     to_signed(895519473, 32), to_signed(895405861, 32), to_signed(895292215, 32), to_signed(895178537, 32),
     to_signed(895064826, 32), to_signed(894951082, 32), to_signed(894837305, 32), to_signed(894723495, 32),
     to_signed(894609652, 32), to_signed(894495777, 32), to_signed(894381868, 32), to_signed(894267927, 32),
     to_signed(894153953, 32), to_signed(894039945, 32), to_signed(893925905, 32), to_signed(893811832, 32),
     to_signed(893697727, 32), to_signed(893583588, 32), to_signed(893469417, 32), to_signed(893355212, 32),
     to_signed(893240975, 32), to_signed(893126705, 32), to_signed(893012402, 32), to_signed(892898067, 32),
     to_signed(892783698, 32), to_signed(892669297, 32), to_signed(892554863, 32), to_signed(892440396, 32),
     to_signed(892325896, 32), to_signed(892211363, 32), to_signed(892096798, 32), to_signed(891982200, 32),
     to_signed(891867569, 32), to_signed(891752905, 32), to_signed(891638208, 32), to_signed(891523479, 32),
     to_signed(891408717, 32), to_signed(891293922, 32), to_signed(891179094, 32), to_signed(891064234, 32),
     to_signed(890949341, 32), to_signed(890834415, 32), to_signed(890719456, 32), to_signed(890604465, 32),
     to_signed(890489440, 32), to_signed(890374383, 32), to_signed(890259294, 32), to_signed(890144171, 32),
     to_signed(890029016, 32), to_signed(889913828, 32), to_signed(889798608, 32), to_signed(889683354, 32),
     to_signed(889568068, 32), to_signed(889452750, 32), to_signed(889337398, 32), to_signed(889222014, 32),
     to_signed(889106597, 32), to_signed(888991148, 32), to_signed(888875666, 32), to_signed(888760151, 32),
     to_signed(888644603, 32), to_signed(888529023, 32), to_signed(888413410, 32), to_signed(888297764, 32),
     to_signed(888182086, 32), to_signed(888066375, 32), to_signed(887950632, 32), to_signed(887834856, 32),
     to_signed(887719047, 32), to_signed(887603205, 32), to_signed(887487331, 32), to_signed(887371425, 32),
     to_signed(887255485, 32), to_signed(887139513, 32), to_signed(887023509, 32), to_signed(886907471, 32),
     to_signed(886791402, 32), to_signed(886675299, 32), to_signed(886559164, 32), to_signed(886442997, 32),
     to_signed(886326796, 32), to_signed(886210564, 32), to_signed(886094298, 32), to_signed(885978000, 32),
     to_signed(885861670, 32), to_signed(885745307, 32), to_signed(885628911, 32), to_signed(885512483, 32),
     to_signed(885396022, 32), to_signed(885279529, 32), to_signed(885163003, 32), to_signed(885046444, 32),
     to_signed(884929853, 32), to_signed(884813230, 32), to_signed(884696574, 32), to_signed(884579885, 32),
     to_signed(884463164, 32), to_signed(884346411, 32), to_signed(884229624, 32), to_signed(884112806, 32),
     to_signed(883995955, 32), to_signed(883879071, 32), to_signed(883762155, 32), to_signed(883645206, 32),
     to_signed(883528225, 32), to_signed(883411212, 32), to_signed(883294165, 32), to_signed(883177087, 32),
     to_signed(883059976, 32), to_signed(882942832, 32), to_signed(882825656, 32), to_signed(882708448, 32),
     to_signed(882591207, 32), to_signed(882473934, 32), to_signed(882356628, 32), to_signed(882239290, 32),
     to_signed(882121919, 32), to_signed(882004516, 32), to_signed(881887080, 32), to_signed(881769613, 32),
     to_signed(881652112, 32), to_signed(881534579, 32), to_signed(881417014, 32), to_signed(881299417, 32),
     to_signed(881181787, 32), to_signed(881064124, 32), to_signed(880946429, 32), to_signed(880828702, 32),
     to_signed(880710943, 32), to_signed(880593151, 32), to_signed(880475326, 32), to_signed(880357470, 32),
     to_signed(880239581, 32), to_signed(880121659, 32), to_signed(880003705, 32), to_signed(879885719, 32),
     to_signed(879767701, 32), to_signed(879649650, 32), to_signed(879531567, 32), to_signed(879413451, 32),
     to_signed(879295303, 32), to_signed(879177123, 32), to_signed(879058911, 32), to_signed(878940666, 32),
     to_signed(878822389, 32), to_signed(878704079, 32), to_signed(878585737, 32), to_signed(878467363, 32),
     to_signed(878348957, 32), to_signed(878230518, 32), to_signed(878112047, 32), to_signed(877993544, 32),
     to_signed(877875009, 32), to_signed(877756441, 32), to_signed(877637841, 32), to_signed(877519208, 32),
     to_signed(877400544, 32), to_signed(877281847, 32), to_signed(877163118, 32), to_signed(877044356, 32),
     to_signed(876925563, 32), to_signed(876806737, 32), to_signed(876687879, 32), to_signed(876568988, 32),
     to_signed(876450066, 32), to_signed(876331111, 32), to_signed(876212124, 32), to_signed(876093105, 32),
     to_signed(875974054, 32), to_signed(875854970, 32), to_signed(875735854, 32), to_signed(875616706, 32),
     to_signed(875497526, 32), to_signed(875378313, 32), to_signed(875259069, 32), to_signed(875139792, 32),
     to_signed(875020483, 32), to_signed(874901142, 32), to_signed(874781769, 32), to_signed(874662363, 32),
     to_signed(874542925, 32), to_signed(874423456, 32), to_signed(874303954, 32), to_signed(874184420, 32),
     to_signed(874064853, 32), to_signed(873945255, 32), to_signed(873825625, 32), to_signed(873705962, 32),
     to_signed(873586267, 32), to_signed(873466540, 32), to_signed(873346781, 32), to_signed(873226990, 32),
     to_signed(873107167, 32), to_signed(872987312, 32), to_signed(872867424, 32), to_signed(872747505, 32),
     to_signed(872627553, 32), to_signed(872507570, 32), to_signed(872387554, 32), to_signed(872267506, 32),
     to_signed(872147426, 32), to_signed(872027314, 32), to_signed(871907170, 32), to_signed(871786994, 32),
     to_signed(871666786, 32), to_signed(871546546, 32), to_signed(871426274, 32), to_signed(871305970, 32),
     to_signed(871185633, 32), to_signed(871065265, 32), to_signed(870944865, 32), to_signed(870824432, 32),
     to_signed(870703968, 32), to_signed(870583472, 32), to_signed(870462943, 32), to_signed(870342383, 32),
     to_signed(870221790, 32), to_signed(870101166, 32), to_signed(869980510, 32), to_signed(869859821, 32),
     to_signed(869739101, 32), to_signed(869618348, 32), to_signed(869497564, 32), to_signed(869376748, 32),
     to_signed(869255900, 32), to_signed(869135019, 32), to_signed(869014107, 32), to_signed(868893163, 32),
     to_signed(868772187, 32), to_signed(868651179, 32), to_signed(868530139, 32), to_signed(868409067, 32),
     to_signed(868287963, 32), to_signed(868166828, 32), to_signed(868045660, 32), to_signed(867924460, 32),
     to_signed(867803229, 32), to_signed(867681966, 32), to_signed(867560670, 32), to_signed(867439343, 32),
     to_signed(867317984, 32), to_signed(867196593, 32), to_signed(867075170, 32), to_signed(866953716, 32),
     to_signed(866832229, 32), to_signed(866710710, 32), to_signed(866589160, 32), to_signed(866467578, 32),
     to_signed(866345964, 32), to_signed(866224318, 32), to_signed(866102640, 32), to_signed(865980931, 32),
     to_signed(865859189, 32), to_signed(865737416, 32), to_signed(865615611, 32), to_signed(865493774, 32),
     to_signed(865371905, 32), to_signed(865250004, 32), to_signed(865128072, 32), to_signed(865006108, 32),
     to_signed(864884112, 32), to_signed(864762084, 32), to_signed(864640024, 32), to_signed(864517933, 32),
     to_signed(864395810, 32), to_signed(864273655, 32), to_signed(864151468, 32), to_signed(864029250, 32),
     to_signed(863906999, 32), to_signed(863784717, 32), to_signed(863662404, 32), to_signed(863540058, 32),
     to_signed(863417681, 32), to_signed(863295272, 32), to_signed(863172831, 32), to_signed(863050358, 32),
     to_signed(862927854, 32), to_signed(862805318, 32), to_signed(862682750, 32), to_signed(862560151, 32),
     to_signed(862437520, 32), to_signed(862314857, 32), to_signed(862192163, 32), to_signed(862069436, 32),
     to_signed(861946678, 32), to_signed(861823889, 32), to_signed(861701067, 32), to_signed(861578214, 32),
     to_signed(861455330, 32), to_signed(861332413, 32), to_signed(861209465, 32), to_signed(861086486, 32),
     to_signed(860963474, 32), to_signed(860840431, 32), to_signed(860717357, 32), to_signed(860594250, 32),
     to_signed(860471112, 32), to_signed(860347943, 32), to_signed(860224742, 32), to_signed(860101509, 32),
     to_signed(859978244, 32), to_signed(859854948, 32), to_signed(859731620, 32), to_signed(859608261, 32),
     to_signed(859484870, 32), to_signed(859361448, 32), to_signed(859237994, 32), to_signed(859114508, 32),
     to_signed(858990991, 32), to_signed(858867442, 32), to_signed(858743861, 32), to_signed(858620249, 32),
     to_signed(858496606, 32), to_signed(858372931, 32), to_signed(858249224, 32), to_signed(858125486, 32),
     to_signed(858001716, 32), to_signed(857877914, 32), to_signed(857754081, 32), to_signed(857630217, 32),
     to_signed(857506321, 32), to_signed(857382394, 32), to_signed(857258434, 32), to_signed(857134444, 32),
     to_signed(857010422, 32), to_signed(856886368, 32), to_signed(856762283, 32), to_signed(856638167, 32),
     to_signed(856514019, 32), to_signed(856389839, 32), to_signed(856265628, 32), to_signed(856141385, 32),
     to_signed(856017111, 32), to_signed(855892806, 32), to_signed(855768469, 32), to_signed(855644100, 32),
     to_signed(855519701, 32), to_signed(855395269, 32), to_signed(855270806, 32), to_signed(855146312, 32),
     to_signed(855021787, 32), to_signed(854897229, 32), to_signed(854772641, 32), to_signed(854648021, 32),
     to_signed(854523370, 32), to_signed(854398687, 32), to_signed(854273973, 32), to_signed(854149227, 32),
     to_signed(854024450, 32), to_signed(853899641, 32), to_signed(853774802, 32), to_signed(853649930, 32),
     to_signed(853525028, 32), to_signed(853400094, 32), to_signed(853275128, 32), to_signed(853150132, 32),
     to_signed(853025104, 32), to_signed(852900044, 32), to_signed(852774953, 32), to_signed(852649831, 32),
     to_signed(852524677, 32), to_signed(852399493, 32), to_signed(852274276, 32), to_signed(852149029, 32),
     to_signed(852023750, 32), to_signed(851898440, 32), to_signed(851773098, 32), to_signed(851647725, 32),
     to_signed(851522321, 32), to_signed(851396886, 32), to_signed(851271419, 32), to_signed(851145921, 32),
     to_signed(851020391, 32), to_signed(850894831, 32), to_signed(850769239, 32), to_signed(850643616, 32),
     to_signed(850517961, 32), to_signed(850392275, 32), to_signed(850266558, 32), to_signed(850140810, 32),
     to_signed(850015030, 32), to_signed(849889220, 32), to_signed(849763378, 32), to_signed(849637504, 32),
     to_signed(849511600, 32), to_signed(849385664, 32), to_signed(849259697, 32), to_signed(849133699, 32),
     to_signed(849007669, 32), to_signed(848881609, 32), to_signed(848755517, 32), to_signed(848629394, 32),
     to_signed(848503239, 32), to_signed(848377054, 32), to_signed(848250837, 32), to_signed(848124589, 32),
     to_signed(847998310, 32), to_signed(847872000, 32), to_signed(847745659, 32), to_signed(847619286, 32),
     to_signed(847492882, 32), to_signed(847366447, 32), to_signed(847239981, 32), to_signed(847113484, 32),
     to_signed(846986956, 32), to_signed(846860396, 32), to_signed(846733806, 32), to_signed(846607184, 32),
     to_signed(846480531, 32), to_signed(846353847, 32), to_signed(846227132, 32), to_signed(846100386, 32),
     to_signed(845973608, 32), to_signed(845846800, 32), to_signed(845719960, 32), to_signed(845593090, 32),
     to_signed(845466188, 32), to_signed(845339255, 32), to_signed(845212291, 32), to_signed(845085296, 32),
     to_signed(844958270, 32), to_signed(844831213, 32), to_signed(844704125, 32), to_signed(844577006, 32),
     to_signed(844449856, 32), to_signed(844322674, 32), to_signed(844195462, 32), to_signed(844068218, 32),
     to_signed(843940944, 32), to_signed(843813638, 32), to_signed(843686302, 32), to_signed(843558934, 32),
     to_signed(843431536, 32), to_signed(843304106, 32), to_signed(843176646, 32), to_signed(843049154, 32),
     to_signed(842921632, 32), to_signed(842794078, 32), to_signed(842666494, 32), to_signed(842538878, 32),
     to_signed(842411232, 32), to_signed(842283554, 32), to_signed(842155846, 32), to_signed(842028106, 32),
     to_signed(841900336, 32), to_signed(841772535, 32), to_signed(841644702, 32), to_signed(841516839, 32),
     to_signed(841388945, 32), to_signed(841261020, 32), to_signed(841133064, 32), to_signed(841005077, 32),
     to_signed(840877059, 32), to_signed(840749010, 32), to_signed(840620931, 32), to_signed(840492820, 32),
     to_signed(840364679, 32), to_signed(840236506, 32), to_signed(840108303, 32), to_signed(839980069, 32),
     to_signed(839851804, 32), to_signed(839723508, 32), to_signed(839595181, 32), to_signed(839466823, 32),
     to_signed(839338435, 32), to_signed(839210015, 32), to_signed(839081565, 32), to_signed(838953084, 32),
     to_signed(838824572, 32), to_signed(838696029, 32), to_signed(838567456, 32), to_signed(838438851, 32),
     to_signed(838310216, 32), to_signed(838181550, 32), to_signed(838052853, 32), to_signed(837924125, 32),
     to_signed(837795367, 32), to_signed(837666577, 32), to_signed(837537757, 32), to_signed(837408906, 32),
     to_signed(837280024, 32), to_signed(837151112, 32), to_signed(837022168, 32), to_signed(836893194, 32),
     to_signed(836764190, 32), to_signed(836635154, 32), to_signed(836506088, 32), to_signed(836376990, 32),
     to_signed(836247863, 32), to_signed(836118704, 32), to_signed(835989515, 32), to_signed(835860294, 32),
     to_signed(835731044, 32), to_signed(835601762, 32), to_signed(835472450, 32), to_signed(835343107, 32),
     to_signed(835213733, 32), to_signed(835084329, 32), to_signed(834954893, 32), to_signed(834825428, 32),
     to_signed(834695931, 32), to_signed(834566404, 32), to_signed(834436846, 32), to_signed(834307257, 32),
     to_signed(834177638, 32), to_signed(834047988, 32), to_signed(833918308, 32), to_signed(833788596, 32),
     to_signed(833658855, 32), to_signed(833529082, 32), to_signed(833399279, 32), to_signed(833269445, 32),
     to_signed(833139580, 32), to_signed(833009685, 32), to_signed(832879760, 32), to_signed(832749803, 32),
     to_signed(832619816, 32), to_signed(832489799, 32), to_signed(832359750, 32), to_signed(832229672, 32),
     to_signed(832099562, 32), to_signed(831969422, 32), to_signed(831839252, 32), to_signed(831709050, 32),
     to_signed(831578819, 32), to_signed(831448556, 32), to_signed(831318263, 32), to_signed(831187940, 32),
     to_signed(831057586, 32), to_signed(830927201, 32), to_signed(830796786, 32), to_signed(830666341, 32),
     to_signed(830535864, 32), to_signed(830405358, 32), to_signed(830274820, 32), to_signed(830144252, 32),
     to_signed(830013654, 32), to_signed(829883025, 32), to_signed(829752366, 32), to_signed(829621676, 32),
     to_signed(829490956, 32), to_signed(829360205, 32), to_signed(829229423, 32), to_signed(829098612, 32),
     to_signed(828967769, 32), to_signed(828836896, 32), to_signed(828705993, 32), to_signed(828575059, 32),
     to_signed(828444095, 32), to_signed(828313100, 32), to_signed(828182075, 32), to_signed(828051020, 32),
     to_signed(827919934, 32), to_signed(827788817, 32), to_signed(827657670, 32), to_signed(827526493, 32),
     to_signed(827395285, 32), to_signed(827264047, 32), to_signed(827132778, 32), to_signed(827001479, 32),
     to_signed(826870150, 32), to_signed(826738790, 32), to_signed(826607400, 32), to_signed(826475979, 32),
     to_signed(826344528, 32), to_signed(826213047, 32), to_signed(826081535, 32), to_signed(825949993, 32),
     to_signed(825818421, 32), to_signed(825686818, 32), to_signed(825555185, 32), to_signed(825423521, 32),
     to_signed(825291827, 32), to_signed(825160103, 32), to_signed(825028348, 32), to_signed(824896563, 32),
     to_signed(824764748, 32), to_signed(824632902, 32), to_signed(824501026, 32), to_signed(824369120, 32),
     to_signed(824237184, 32), to_signed(824105217, 32), to_signed(823973220, 32), to_signed(823841192, 32),
     to_signed(823709135, 32), to_signed(823577047, 32), to_signed(823444928, 32), to_signed(823312780, 32),
     to_signed(823180601, 32), to_signed(823048392, 32), to_signed(822916152, 32), to_signed(822783883, 32),
     to_signed(822651583, 32), to_signed(822519253, 32), to_signed(822386892, 32), to_signed(822254502, 32),
     to_signed(822122081, 32), to_signed(821989630, 32), to_signed(821857149, 32), to_signed(821724637, 32),
     to_signed(821592095, 32), to_signed(821459524, 32), to_signed(821326921, 32), to_signed(821194289, 32),
     to_signed(821061627, 32), to_signed(820928934, 32), to_signed(820796211, 32), to_signed(820663458, 32),
     to_signed(820530675, 32), to_signed(820397861, 32), to_signed(820265018, 32), to_signed(820132144, 32),
     to_signed(819999240, 32), to_signed(819866306, 32), to_signed(819733342, 32), to_signed(819600348, 32),
     to_signed(819467323, 32), to_signed(819334269, 32), to_signed(819201184, 32), to_signed(819068069, 32),
     to_signed(818934924, 32), to_signed(818801749, 32), to_signed(818668544, 32), to_signed(818535309, 32),
     to_signed(818402043, 32), to_signed(818268748, 32), to_signed(818135422, 32), to_signed(818002067, 32),
     to_signed(817868681, 32), to_signed(817735265, 32), to_signed(817601820, 32), to_signed(817468344, 32),
     to_signed(817334838, 32), to_signed(817201302, 32), to_signed(817067736, 32), to_signed(816934140, 32),
     to_signed(816800514, 32), to_signed(816666858, 32), to_signed(816533171, 32), to_signed(816399455, 32),
     to_signed(816265709, 32), to_signed(816131933, 32), to_signed(815998127, 32), to_signed(815864290, 32),
     to_signed(815730424, 32), to_signed(815596528, 32), to_signed(815462602, 32), to_signed(815328646, 32),
     to_signed(815194659, 32), to_signed(815060643, 32), to_signed(814926597, 32), to_signed(814792521, 32),
     to_signed(814658415, 32), to_signed(814524279, 32), to_signed(814390113, 32), to_signed(814255917, 32),
     to_signed(814121692, 32), to_signed(813987436, 32), to_signed(813853150, 32), to_signed(813718835, 32),
     to_signed(813584489, 32), to_signed(813450114, 32), to_signed(813315708, 32), to_signed(813181273, 32),
     to_signed(813046808, 32), to_signed(812912313, 32), to_signed(812777788, 32), to_signed(812643233, 32),
     to_signed(812508649, 32), to_signed(812374034, 32), to_signed(812239390, 32), to_signed(812104715, 32),
     to_signed(811970011, 32), to_signed(811835277, 32), to_signed(811700513, 32), to_signed(811565720, 32),
     to_signed(811430896, 32), to_signed(811296043, 32), to_signed(811161160, 32), to_signed(811026247, 32),
     to_signed(810891304, 32), to_signed(810756331, 32), to_signed(810621329, 32), to_signed(810486297, 32),
     to_signed(810351235, 32), to_signed(810216143, 32), to_signed(810081021, 32), to_signed(809945870, 32),
     to_signed(809810688, 32), to_signed(809675477, 32), to_signed(809540237, 32), to_signed(809404966, 32),
     to_signed(809269666, 32), to_signed(809134336, 32), to_signed(808998976, 32), to_signed(808863587, 32),
     to_signed(808728167, 32), to_signed(808592718, 32), to_signed(808457240, 32), to_signed(808321731, 32),
     to_signed(808186193, 32), to_signed(808050625, 32), to_signed(807915028, 32), to_signed(807779400, 32),
     to_signed(807643743, 32), to_signed(807508057, 32), to_signed(807372340, 32), to_signed(807236594, 32),
     to_signed(807100819, 32), to_signed(806965013, 32), to_signed(806829178, 32), to_signed(806693313, 32),
     to_signed(806557419, 32), to_signed(806421495, 32), to_signed(806285541, 32), to_signed(806149558, 32),
     to_signed(806013545, 32), to_signed(805877502, 32), to_signed(805741430, 32), to_signed(805605328, 32),
     to_signed(805469196, 32), to_signed(805333035, 32), to_signed(805196845, 32), to_signed(805060624, 32),
     to_signed(804924374, 32), to_signed(804788095, 32), to_signed(804651786, 32), to_signed(804515447, 32),
     to_signed(804379079, 32), to_signed(804242681, 32), to_signed(804106253, 32), to_signed(803969796, 32),
     to_signed(803833310, 32), to_signed(803696794, 32), to_signed(803560248, 32), to_signed(803423673, 32),
     to_signed(803287068, 32), to_signed(803150434, 32), to_signed(803013770, 32), to_signed(802877077, 32),
     to_signed(802740354, 32), to_signed(802603602, 32), to_signed(802466820, 32), to_signed(802330008, 32),
     to_signed(802193167, 32), to_signed(802056297, 32), to_signed(801919397, 32), to_signed(801782468, 32),
     to_signed(801645509, 32), to_signed(801508521, 32), to_signed(801371503, 32), to_signed(801234456, 32),
     to_signed(801097379, 32), to_signed(800960273, 32), to_signed(800823137, 32), to_signed(800685972, 32),
     to_signed(800548778, 32), to_signed(800411554, 32), to_signed(800274300, 32), to_signed(800137018, 32),
     to_signed(799999706, 32), to_signed(799862364, 32), to_signed(799724993, 32), to_signed(799587593, 32),
     to_signed(799450163, 32), to_signed(799312704, 32), to_signed(799175215, 32), to_signed(799037697, 32),
     to_signed(798900150, 32), to_signed(798762573, 32), to_signed(798624967, 32), to_signed(798487331, 32),
     to_signed(798349667, 32), to_signed(798211972, 32), to_signed(798074249, 32), to_signed(797936496, 32),
     to_signed(797798714, 32), to_signed(797660902, 32), to_signed(797523061, 32), to_signed(797385191, 32),
     to_signed(797247292, 32), to_signed(797109363, 32), to_signed(796971405, 32), to_signed(796833417, 32),
     to_signed(796695401, 32), to_signed(796557355, 32), to_signed(796419279, 32), to_signed(796281175, 32),
     to_signed(796143041, 32), to_signed(796004878, 32), to_signed(795866685, 32), to_signed(795728464, 32),
     to_signed(795590213, 32), to_signed(795451933, 32), to_signed(795313623, 32), to_signed(795175285, 32),
     to_signed(795036917, 32), to_signed(794898520, 32), to_signed(794760093, 32), to_signed(794621638, 32),
     to_signed(794483153, 32), to_signed(794344639, 32), to_signed(794206096, 32), to_signed(794067523, 32),
     to_signed(793928922, 32), to_signed(793790291, 32), to_signed(793651631, 32), to_signed(793512942, 32),
     to_signed(793374223, 32), to_signed(793235476, 32), to_signed(793096699, 32), to_signed(792957894, 32),
     to_signed(792819059, 32), to_signed(792680194, 32), to_signed(792541301, 32), to_signed(792402379, 32),
     to_signed(792263427, 32), to_signed(792124447, 32), to_signed(791985437, 32), to_signed(791846398, 32),
     to_signed(791707330, 32), to_signed(791568233, 32), to_signed(791429106, 32), to_signed(791289951, 32),
     to_signed(791150767, 32), to_signed(791011553, 32), to_signed(790872310, 32), to_signed(790733039, 32),
     to_signed(790593738, 32), to_signed(790454408, 32), to_signed(790315049, 32), to_signed(790175661, 32),
     to_signed(790036244, 32), to_signed(789896798, 32), to_signed(789757323, 32), to_signed(789617819, 32),
     to_signed(789478286, 32), to_signed(789338724, 32), to_signed(789199133, 32), to_signed(789059512, 32),
     to_signed(788919863, 32), to_signed(788780185, 32), to_signed(788640478, 32), to_signed(788500741, 32),
     to_signed(788360976, 32), to_signed(788221182, 32), to_signed(788081359, 32), to_signed(787941507, 32),
     to_signed(787801625, 32), to_signed(787661715, 32), to_signed(787521776, 32), to_signed(787381808, 32),
     to_signed(787241811, 32), to_signed(787101785, 32), to_signed(786961731, 32), to_signed(786821647, 32),
     to_signed(786681534, 32), to_signed(786541392, 32), to_signed(786401222, 32), to_signed(786261022, 32),
     to_signed(786120794, 32), to_signed(785980537, 32), to_signed(785840250, 32), to_signed(785699935, 32),
     to_signed(785559591, 32), to_signed(785419219, 32), to_signed(785278817, 32), to_signed(785138386, 32),
     to_signed(784997927, 32), to_signed(784857438, 32), to_signed(784716921, 32), to_signed(784576375, 32),
     to_signed(784435800, 32), to_signed(784295197, 32), to_signed(784154564, 32), to_signed(784013903, 32),
     to_signed(783873212, 32), to_signed(783732493, 32), to_signed(783591746, 32), to_signed(783450969, 32),
     to_signed(783310163, 32), to_signed(783169329, 32), to_signed(783028466, 32), to_signed(782887574, 32),
     to_signed(782746654, 32), to_signed(782605704, 32), to_signed(782464726, 32), to_signed(782323719, 32),
     to_signed(782182683, 32), to_signed(782041619, 32), to_signed(781900526, 32), to_signed(781759404, 32),
     to_signed(781618253, 32), to_signed(781477073, 32), to_signed(781335865, 32), to_signed(781194628, 32),
     to_signed(781053363, 32), to_signed(780912068, 32), to_signed(780770745, 32), to_signed(780629393, 32),
     to_signed(780488013, 32), to_signed(780346604, 32), to_signed(780205166, 32), to_signed(780063699, 32),
     to_signed(779922204, 32), to_signed(779780680, 32), to_signed(779639128, 32), to_signed(779497546, 32),
     to_signed(779355936, 32), to_signed(779214298, 32), to_signed(779072631, 32), to_signed(778930935, 32),
     to_signed(778789210, 32), to_signed(778647457, 32), to_signed(778505675, 32), to_signed(778363865, 32),
     to_signed(778222026, 32), to_signed(778080158, 32), to_signed(777938262, 32), to_signed(777796337, 32),
     to_signed(777654384, 32), to_signed(777512402, 32), to_signed(777370391, 32), to_signed(777228352, 32),
     to_signed(777086284, 32), to_signed(776944188, 32), to_signed(776802063, 32), to_signed(776659910, 32),
     to_signed(776517728, 32), to_signed(776375517, 32), to_signed(776233278, 32), to_signed(776091010, 32),
     to_signed(775948714, 32), to_signed(775806389, 32), to_signed(775664036, 32), to_signed(775521654, 32),
     to_signed(775379244, 32), to_signed(775236805, 32), to_signed(775094338, 32), to_signed(774951842, 32),
     to_signed(774809318, 32), to_signed(774666765, 32), to_signed(774524184, 32), to_signed(774381574, 32),
     to_signed(774238936, 32), to_signed(774096269, 32), to_signed(773953574, 32), to_signed(773810851, 32),
     to_signed(773668099, 32), to_signed(773525318, 32), to_signed(773382509, 32), to_signed(773239672, 32),
     to_signed(773096806, 32), to_signed(772953912, 32), to_signed(772810989, 32), to_signed(772668038, 32),
     to_signed(772525059, 32), to_signed(772382051, 32), to_signed(772239015, 32), to_signed(772095950, 32),
     to_signed(771952857, 32), to_signed(771809736, 32), to_signed(771666586, 32), to_signed(771523408, 32),
     to_signed(771380201, 32), to_signed(771236966, 32), to_signed(771093703, 32), to_signed(770950412, 32),
     to_signed(770807092, 32), to_signed(770663743, 32), to_signed(770520367, 32), to_signed(770376962, 32),
     to_signed(770233528, 32), to_signed(770090067, 32), to_signed(769946577, 32), to_signed(769803059, 32),
     to_signed(769659512, 32), to_signed(769515937, 32), to_signed(769372334, 32), to_signed(769228703, 32),
     to_signed(769085043, 32), to_signed(768941355, 32), to_signed(768797639, 32), to_signed(768653895, 32),
     to_signed(768510122, 32), to_signed(768366321, 32), to_signed(768222492, 32), to_signed(768078634, 32),
     to_signed(767934748, 32), to_signed(767790834, 32), to_signed(767646892, 32), to_signed(767502922, 32),
     to_signed(767358923, 32), to_signed(767214896, 32), to_signed(767070841, 32), to_signed(766926758, 32),
     to_signed(766782646, 32), to_signed(766638507, 32), to_signed(766494339, 32), to_signed(766350143, 32),
     to_signed(766205919, 32), to_signed(766061666, 32), to_signed(765917386, 32), to_signed(765773077, 32),
     to_signed(765628740, 32), to_signed(765484375, 32), to_signed(765339982, 32), to_signed(765195561, 32),
     to_signed(765051111, 32), to_signed(764906634, 32), to_signed(764762128, 32), to_signed(764617594, 32),
     to_signed(764473032, 32), to_signed(764328442, 32), to_signed(764183824, 32), to_signed(764039178, 32),
     to_signed(763894504, 32), to_signed(763749801, 32), to_signed(763605071, 32), to_signed(763460312, 32),
     to_signed(763315525, 32), to_signed(763170711, 32), to_signed(763025868, 32), to_signed(762880997, 32),
     to_signed(762736098, 32), to_signed(762591171, 32), to_signed(762446217, 32), to_signed(762301234, 32),
     to_signed(762156223, 32), to_signed(762011184, 32), to_signed(761866116, 32), to_signed(761721021, 32),
     to_signed(761575898, 32), to_signed(761430747, 32), to_signed(761285568, 32), to_signed(761140361, 32),
     to_signed(760995126, 32), to_signed(760849863, 32), to_signed(760704572, 32), to_signed(760559253, 32),
     to_signed(760413906, 32), to_signed(760268531, 32), to_signed(760123129, 32), to_signed(759977698, 32),
     to_signed(759832239, 32), to_signed(759686753, 32), to_signed(759541238, 32), to_signed(759395695, 32));  -- sfix32 [4096]
  CONSTANT Twiddle_im_table_data          : vector_of_signed32(0 TO 4095) := 
    (to_signed(0, 32), to_signed(-205887, 32), to_signed(-411775, 32), to_signed(-617662, 32),
     to_signed(-823550, 32), to_signed(-1029437, 32), to_signed(-1235324, 32), to_signed(-1441211, 32),
     to_signed(-1647099, 32), to_signed(-1852986, 32), to_signed(-2058873, 32), to_signed(-2264760, 32),
     to_signed(-2470647, 32), to_signed(-2676534, 32), to_signed(-2882420, 32), to_signed(-3088307, 32),
     to_signed(-3294193, 32), to_signed(-3500080, 32), to_signed(-3705966, 32), to_signed(-3911852, 32),
     to_signed(-4117738, 32), to_signed(-4323624, 32), to_signed(-4529510, 32), to_signed(-4735395, 32),
     to_signed(-4941281, 32), to_signed(-5147166, 32), to_signed(-5353051, 32), to_signed(-5558935, 32),
     to_signed(-5764820, 32), to_signed(-5970704, 32), to_signed(-6176588, 32), to_signed(-6382472, 32),
     to_signed(-6588356, 32), to_signed(-6794239, 32), to_signed(-7000123, 32), to_signed(-7206005, 32),
     to_signed(-7411888, 32), to_signed(-7617770, 32), to_signed(-7823653, 32), to_signed(-8029534, 32),
     to_signed(-8235416, 32), to_signed(-8441297, 32), to_signed(-8647178, 32), to_signed(-8853059, 32),
     to_signed(-9058939, 32), to_signed(-9264819, 32), to_signed(-9470698, 32), to_signed(-9676578, 32),
     to_signed(-9882456, 32), to_signed(-10088335, 32), to_signed(-10294213, 32), to_signed(-10500091, 32),
     to_signed(-10705968, 32), to_signed(-10911845, 32), to_signed(-11117722, 32), to_signed(-11323598, 32),
     to_signed(-11529474, 32), to_signed(-11735349, 32), to_signed(-11941224, 32), to_signed(-12147098, 32),
     to_signed(-12352972, 32), to_signed(-12558846, 32), to_signed(-12764719, 32), to_signed(-12970592, 32),
     to_signed(-13176464, 32), to_signed(-13382336, 32), to_signed(-13588207, 32), to_signed(-13794077, 32),
     to_signed(-13999948, 32), to_signed(-14205817, 32), to_signed(-14411686, 32), to_signed(-14617555, 32),
     to_signed(-14823423, 32), to_signed(-15029291, 32), to_signed(-15235158, 32), to_signed(-15441024, 32),
     to_signed(-15646890, 32), to_signed(-15852755, 32), to_signed(-16058620, 32), to_signed(-16264484, 32),
     to_signed(-16470347, 32), to_signed(-16676210, 32), to_signed(-16882072, 32), to_signed(-17087934, 32),
     to_signed(-17293795, 32), to_signed(-17499656, 32), to_signed(-17705515, 32), to_signed(-17911374, 32),
     to_signed(-18117233, 32), to_signed(-18323091, 32), to_signed(-18528948, 32), to_signed(-18734804, 32),
     to_signed(-18940660, 32), to_signed(-19146515, 32), to_signed(-19352369, 32), to_signed(-19558223, 32),
     to_signed(-19764076, 32), to_signed(-19969928, 32), to_signed(-20175779, 32), to_signed(-20381630, 32),
     to_signed(-20587480, 32), to_signed(-20793329, 32), to_signed(-20999178, 32), to_signed(-21205025, 32),
     to_signed(-21410872, 32), to_signed(-21616718, 32), to_signed(-21822563, 32), to_signed(-22028408, 32),
     to_signed(-22234252, 32), to_signed(-22440095, 32), to_signed(-22645937, 32), to_signed(-22851778, 32),
     to_signed(-23057618, 32), to_signed(-23263458, 32), to_signed(-23469296, 32), to_signed(-23675134, 32),
     to_signed(-23880971, 32), to_signed(-24086807, 32), to_signed(-24292642, 32), to_signed(-24498476, 32),
     to_signed(-24704310, 32), to_signed(-24910142, 32), to_signed(-25115974, 32), to_signed(-25321804, 32),
     to_signed(-25527634, 32), to_signed(-25733463, 32), to_signed(-25939291, 32), to_signed(-26145118, 32),
     to_signed(-26350943, 32), to_signed(-26556768, 32), to_signed(-26762592, 32), to_signed(-26968415, 32),
     to_signed(-27174237, 32), to_signed(-27380058, 32), to_signed(-27585878, 32), to_signed(-27791697, 32),
     to_signed(-27997515, 32), to_signed(-28203332, 32), to_signed(-28409148, 32), to_signed(-28614963, 32),
     to_signed(-28820776, 32), to_signed(-29026589, 32), to_signed(-29232401, 32), to_signed(-29438211, 32),
     to_signed(-29644021, 32), to_signed(-29849829, 32), to_signed(-30055636, 32), to_signed(-30261443, 32),
     to_signed(-30467248, 32), to_signed(-30673052, 32), to_signed(-30878855, 32), to_signed(-31084656, 32),
     to_signed(-31290457, 32), to_signed(-31496256, 32), to_signed(-31702054, 32), to_signed(-31907851, 32),
     to_signed(-32113647, 32), to_signed(-32319442, 32), to_signed(-32525236, 32), to_signed(-32731028, 32),
     to_signed(-32936819, 32), to_signed(-33142609, 32), to_signed(-33348398, 32), to_signed(-33554185, 32),
     to_signed(-33759971, 32), to_signed(-33965756, 32), to_signed(-34171540, 32), to_signed(-34377323, 32),
     to_signed(-34583104, 32), to_signed(-34788884, 32), to_signed(-34994663, 32), to_signed(-35200440, 32),
     to_signed(-35406216, 32), to_signed(-35611991, 32), to_signed(-35817764, 32), to_signed(-36023537, 32),
     to_signed(-36229307, 32), to_signed(-36435077, 32), to_signed(-36640845, 32), to_signed(-36846612, 32),
     to_signed(-37052377, 32), to_signed(-37258142, 32), to_signed(-37463904, 32), to_signed(-37669666, 32),
     to_signed(-37875426, 32), to_signed(-38081184, 32), to_signed(-38286941, 32), to_signed(-38492697, 32),
     to_signed(-38698452, 32), to_signed(-38904204, 32), to_signed(-39109956, 32), to_signed(-39315706, 32),
     to_signed(-39521455, 32), to_signed(-39727202, 32), to_signed(-39932948, 32), to_signed(-40138692, 32),
     to_signed(-40344435, 32), to_signed(-40550176, 32), to_signed(-40755916, 32), to_signed(-40961654, 32),
     to_signed(-41167391, 32), to_signed(-41373126, 32), to_signed(-41578860, 32), to_signed(-41784592, 32),
     to_signed(-41990323, 32), to_signed(-42196052, 32), to_signed(-42401779, 32), to_signed(-42607506, 32),
     to_signed(-42813230, 32), to_signed(-43018953, 32), to_signed(-43224674, 32), to_signed(-43430394, 32),
     to_signed(-43636112, 32), to_signed(-43841829, 32), to_signed(-44047544, 32), to_signed(-44253257, 32),
     to_signed(-44458968, 32), to_signed(-44664678, 32), to_signed(-44870387, 32), to_signed(-45076094, 32),
     to_signed(-45281799, 32), to_signed(-45487502, 32), to_signed(-45693204, 32), to_signed(-45898904, 32),
     to_signed(-46104602, 32), to_signed(-46310299, 32), to_signed(-46515994, 32), to_signed(-46721687, 32),
     to_signed(-46927379, 32), to_signed(-47133069, 32), to_signed(-47338757, 32), to_signed(-47544443, 32),
     to_signed(-47750128, 32), to_signed(-47955811, 32), to_signed(-48161492, 32), to_signed(-48367171, 32),
     to_signed(-48572848, 32), to_signed(-48778524, 32), to_signed(-48984198, 32), to_signed(-49189870, 32),
     to_signed(-49395541, 32), to_signed(-49601209, 32), to_signed(-49806876, 32), to_signed(-50012541, 32),
     to_signed(-50218204, 32), to_signed(-50423865, 32), to_signed(-50629524, 32), to_signed(-50835182, 32),
     to_signed(-51040837, 32), to_signed(-51246491, 32), to_signed(-51452143, 32), to_signed(-51657793, 32),
     to_signed(-51863441, 32), to_signed(-52069087, 32), to_signed(-52274731, 32), to_signed(-52480374, 32),
     to_signed(-52686014, 32), to_signed(-52891653, 32), to_signed(-53097289, 32), to_signed(-53302924, 32),
     to_signed(-53508556, 32), to_signed(-53714187, 32), to_signed(-53919815, 32), to_signed(-54125442, 32),
     to_signed(-54331067, 32), to_signed(-54536690, 32), to_signed(-54742310, 32), to_signed(-54947929, 32),
     to_signed(-55153545, 32), to_signed(-55359160, 32), to_signed(-55564773, 32), to_signed(-55770383, 32),
     to_signed(-55975992, 32), to_signed(-56181598, 32), to_signed(-56387202, 32), to_signed(-56592805, 32),
     to_signed(-56798405, 32), to_signed(-57004003, 32), to_signed(-57209599, 32), to_signed(-57415193, 32),
     to_signed(-57620785, 32), to_signed(-57826374, 32), to_signed(-58031962, 32), to_signed(-58237547, 32),
     to_signed(-58443131, 32), to_signed(-58648712, 32), to_signed(-58854291, 32), to_signed(-59059868, 32),
     to_signed(-59265442, 32), to_signed(-59471015, 32), to_signed(-59676585, 32), to_signed(-59882153, 32),
     to_signed(-60087719, 32), to_signed(-60293283, 32), to_signed(-60498844, 32), to_signed(-60704403, 32),
     to_signed(-60909960, 32), to_signed(-61115515, 32), to_signed(-61321068, 32), to_signed(-61526618, 32),
     to_signed(-61732166, 32), to_signed(-61937712, 32), to_signed(-62143255, 32), to_signed(-62348796, 32),
     to_signed(-62554335, 32), to_signed(-62759872, 32), to_signed(-62965406, 32), to_signed(-63170938, 32),
     to_signed(-63376468, 32), to_signed(-63581995, 32), to_signed(-63787520, 32), to_signed(-63993042, 32),
     to_signed(-64198563, 32), to_signed(-64404081, 32), to_signed(-64609596, 32), to_signed(-64815109, 32),
     to_signed(-65020620, 32), to_signed(-65226129, 32), to_signed(-65431634, 32), to_signed(-65637138, 32),
     to_signed(-65842639, 32), to_signed(-66048138, 32), to_signed(-66253634, 32), to_signed(-66459128, 32),
     to_signed(-66664620, 32), to_signed(-66870109, 32), to_signed(-67075595, 32), to_signed(-67281079, 32),
     to_signed(-67486561, 32), to_signed(-67692040, 32), to_signed(-67897517, 32), to_signed(-68102991, 32),
     to_signed(-68308462, 32), to_signed(-68513931, 32), to_signed(-68719398, 32), to_signed(-68924862, 32),
     to_signed(-69130324, 32), to_signed(-69335783, 32), to_signed(-69541239, 32), to_signed(-69746693, 32),
     to_signed(-69952144, 32), to_signed(-70157593, 32), to_signed(-70363039, 32), to_signed(-70568483, 32),
     to_signed(-70773924, 32), to_signed(-70979362, 32), to_signed(-71184798, 32), to_signed(-71390231, 32),
     to_signed(-71595661, 32), to_signed(-71801089, 32), to_signed(-72006515, 32), to_signed(-72211937, 32),
     to_signed(-72417357, 32), to_signed(-72622775, 32), to_signed(-72828189, 32), to_signed(-73033601, 32),
     to_signed(-73239010, 32), to_signed(-73444417, 32), to_signed(-73649821, 32), to_signed(-73855222, 32),
     to_signed(-74060620, 32), to_signed(-74266016, 32), to_signed(-74471409, 32), to_signed(-74676799, 32),
     to_signed(-74882187, 32), to_signed(-75087572, 32), to_signed(-75292954, 32), to_signed(-75498333, 32),
     to_signed(-75703709, 32), to_signed(-75909083, 32), to_signed(-76114454, 32), to_signed(-76319822, 32),
     to_signed(-76525187, 32), to_signed(-76730550, 32), to_signed(-76935909, 32), to_signed(-77141266, 32),
     to_signed(-77346620, 32), to_signed(-77551971, 32), to_signed(-77757319, 32), to_signed(-77962665, 32),
     to_signed(-78168007, 32), to_signed(-78373347, 32), to_signed(-78578684, 32), to_signed(-78784018, 32),
     to_signed(-78989349, 32), to_signed(-79194677, 32), to_signed(-79400002, 32), to_signed(-79605324, 32),
     to_signed(-79810644, 32), to_signed(-80015960, 32), to_signed(-80221273, 32), to_signed(-80426584, 32),
     to_signed(-80631892, 32), to_signed(-80837196, 32), to_signed(-81042498, 32), to_signed(-81247796, 32),
     to_signed(-81453092, 32), to_signed(-81658385, 32), to_signed(-81863674, 32), to_signed(-82068961, 32),
     to_signed(-82274245, 32), to_signed(-82479525, 32), to_signed(-82684803, 32), to_signed(-82890077, 32),
     to_signed(-83095349, 32), to_signed(-83300617, 32), to_signed(-83505883, 32), to_signed(-83711145, 32),
     to_signed(-83916404, 32), to_signed(-84121660, 32), to_signed(-84326913, 32), to_signed(-84532163, 32),
     to_signed(-84737410, 32), to_signed(-84942654, 32), to_signed(-85147894, 32), to_signed(-85353132, 32),
     to_signed(-85558366, 32), to_signed(-85763597, 32), to_signed(-85968825, 32), to_signed(-86174050, 32),
     to_signed(-86379272, 32), to_signed(-86584491, 32), to_signed(-86789706, 32), to_signed(-86994918, 32),
     to_signed(-87200127, 32), to_signed(-87405333, 32), to_signed(-87610535, 32), to_signed(-87815735, 32),
     to_signed(-88020931, 32), to_signed(-88226124, 32), to_signed(-88431313, 32), to_signed(-88636499, 32),
     to_signed(-88841683, 32), to_signed(-89046862, 32), to_signed(-89252039, 32), to_signed(-89457212, 32),
     to_signed(-89662382, 32), to_signed(-89867549, 32), to_signed(-90072712, 32), to_signed(-90277872, 32),
     to_signed(-90483029, 32), to_signed(-90688182, 32), to_signed(-90893333, 32), to_signed(-91098479, 32),
     to_signed(-91303623, 32), to_signed(-91508763, 32), to_signed(-91713899, 32), to_signed(-91919033, 32),
     to_signed(-92124163, 32), to_signed(-92329289, 32), to_signed(-92534412, 32), to_signed(-92739532, 32),
     to_signed(-92944648, 32), to_signed(-93149761, 32), to_signed(-93354871, 32), to_signed(-93559977, 32),
     to_signed(-93765079, 32), to_signed(-93970179, 32), to_signed(-94175274, 32), to_signed(-94380367, 32),
     to_signed(-94585455, 32), to_signed(-94790541, 32), to_signed(-94995622, 32), to_signed(-95200701, 32),
     to_signed(-95405776, 32), to_signed(-95610847, 32), to_signed(-95815915, 32), to_signed(-96020979, 32),
     to_signed(-96226040, 32), to_signed(-96431097, 32), to_signed(-96636151, 32), to_signed(-96841201, 32),
     to_signed(-97046247, 32), to_signed(-97251290, 32), to_signed(-97456330, 32), to_signed(-97661365, 32),
     to_signed(-97866398, 32), to_signed(-98071426, 32), to_signed(-98276451, 32), to_signed(-98481473, 32),
     to_signed(-98686491, 32), to_signed(-98891505, 32), to_signed(-99096515, 32), to_signed(-99301522, 32),
     to_signed(-99506525, 32), to_signed(-99711525, 32), to_signed(-99916521, 32), to_signed(-100121513, 32),
     to_signed(-100326502, 32), to_signed(-100531487, 32), to_signed(-100736468, 32), to_signed(-100941445, 32),
     to_signed(-101146419, 32), to_signed(-101351389, 32), to_signed(-101556355, 32), to_signed(-101761318, 32),
     to_signed(-101966277, 32), to_signed(-102171232, 32), to_signed(-102376183, 32), to_signed(-102581131, 32),
     to_signed(-102786074, 32), to_signed(-102991014, 32), to_signed(-103195951, 32), to_signed(-103400883, 32),
     to_signed(-103605812, 32), to_signed(-103810737, 32), to_signed(-104015658, 32), to_signed(-104220575, 32),
     to_signed(-104425488, 32), to_signed(-104630398, 32), to_signed(-104835303, 32), to_signed(-105040205, 32),
     to_signed(-105245103, 32), to_signed(-105449997, 32), to_signed(-105654887, 32), to_signed(-105859774, 32),
     to_signed(-106064656, 32), to_signed(-106269535, 32), to_signed(-106474409, 32), to_signed(-106679280, 32),
     to_signed(-106884147, 32), to_signed(-107089010, 32), to_signed(-107293868, 32), to_signed(-107498723, 32),
     to_signed(-107703574, 32), to_signed(-107908421, 32), to_signed(-108113265, 32), to_signed(-108318104, 32),
     to_signed(-108522939, 32), to_signed(-108727770, 32), to_signed(-108932597, 32), to_signed(-109137420, 32),
     to_signed(-109342239, 32), to_signed(-109547054, 32), to_signed(-109751866, 32), to_signed(-109956673, 32),
     to_signed(-110161476, 32), to_signed(-110366274, 32), to_signed(-110571069, 32), to_signed(-110775860, 32),
     to_signed(-110980647, 32), to_signed(-111185430, 32), to_signed(-111390208, 32), to_signed(-111594983, 32),
     to_signed(-111799753, 32), to_signed(-112004519, 32), to_signed(-112209281, 32), to_signed(-112414040, 32),
     to_signed(-112618793, 32), to_signed(-112823543, 32), to_signed(-113028289, 32), to_signed(-113233030, 32),
     to_signed(-113437768, 32), to_signed(-113642501, 32), to_signed(-113847230, 32), to_signed(-114051954, 32),
     to_signed(-114256675, 32), to_signed(-114461391, 32), to_signed(-114666103, 32), to_signed(-114870811, 32),
     to_signed(-115075515, 32), to_signed(-115280215, 32), to_signed(-115484910, 32), to_signed(-115689601, 32),
     to_signed(-115894288, 32), to_signed(-116098970, 32), to_signed(-116303648, 32), to_signed(-116508322, 32),
     to_signed(-116712992, 32), to_signed(-116917657, 32), to_signed(-117122318, 32), to_signed(-117326975, 32),
     to_signed(-117531627, 32), to_signed(-117736276, 32), to_signed(-117940919, 32), to_signed(-118145559, 32),
     to_signed(-118350194, 32), to_signed(-118554825, 32), to_signed(-118759451, 32), to_signed(-118964073, 32),
     to_signed(-119168691, 32), to_signed(-119373304, 32), to_signed(-119577913, 32), to_signed(-119782517, 32),
     to_signed(-119987118, 32), to_signed(-120191713, 32), to_signed(-120396304, 32), to_signed(-120600891, 32),
     to_signed(-120805474, 32), to_signed(-121010052, 32), to_signed(-121214625, 32), to_signed(-121419194, 32),
     to_signed(-121623759, 32), to_signed(-121828319, 32), to_signed(-122032875, 32), to_signed(-122237426, 32),
     to_signed(-122441972, 32), to_signed(-122646515, 32), to_signed(-122851052, 32), to_signed(-123055585, 32),
     to_signed(-123260114, 32), to_signed(-123464638, 32), to_signed(-123669157, 32), to_signed(-123873672, 32),
     to_signed(-124078183, 32), to_signed(-124282689, 32), to_signed(-124487190, 32), to_signed(-124691687, 32),
     to_signed(-124896179, 32), to_signed(-125100666, 32), to_signed(-125305149, 32), to_signed(-125509628, 32),
     to_signed(-125714101, 32), to_signed(-125918571, 32), to_signed(-126123035, 32), to_signed(-126327495, 32),
     to_signed(-126531950, 32), to_signed(-126736401, 32), to_signed(-126940846, 32), to_signed(-127145288, 32),
     to_signed(-127349724, 32), to_signed(-127554156, 32), to_signed(-127758583, 32), to_signed(-127963006, 32),
     to_signed(-128167423, 32), to_signed(-128371837, 32), to_signed(-128576245, 32), to_signed(-128780648, 32),
     to_signed(-128985047, 32), to_signed(-129189441, 32), to_signed(-129393831, 32), to_signed(-129598215, 32),
     to_signed(-129802595, 32), to_signed(-130006970, 32), to_signed(-130211341, 32), to_signed(-130415706, 32),
     to_signed(-130620067, 32), to_signed(-130824423, 32), to_signed(-131028774, 32), to_signed(-131233120, 32),
     to_signed(-131437462, 32), to_signed(-131641798, 32), to_signed(-131846130, 32), to_signed(-132050457, 32),
     to_signed(-132254779, 32), to_signed(-132459096, 32), to_signed(-132663409, 32), to_signed(-132867716, 32),
     to_signed(-133072019, 32), to_signed(-133276316, 32), to_signed(-133480609, 32), to_signed(-133684897, 32),
     to_signed(-133889180, 32), to_signed(-134093458, 32), to_signed(-134297731, 32), to_signed(-134501999, 32),
     to_signed(-134706263, 32), to_signed(-134910521, 32), to_signed(-135114774, 32), to_signed(-135319023, 32),
     to_signed(-135523266, 32), to_signed(-135727504, 32), to_signed(-135931738, 32), to_signed(-136135966, 32),
     to_signed(-136340190, 32), to_signed(-136544408, 32), to_signed(-136748621, 32), to_signed(-136952830, 32),
     to_signed(-137157033, 32), to_signed(-137361231, 32), to_signed(-137565425, 32), to_signed(-137769613, 32),
     to_signed(-137973796, 32), to_signed(-138177974, 32), to_signed(-138382147, 32), to_signed(-138586315, 32),
     to_signed(-138790477, 32), to_signed(-138994635, 32), to_signed(-139198788, 32), to_signed(-139402935, 32),
     to_signed(-139607077, 32), to_signed(-139811215, 32), to_signed(-140015347, 32), to_signed(-140219473, 32),
     to_signed(-140423595, 32), to_signed(-140627712, 32), to_signed(-140831823, 32), to_signed(-141035929, 32),
     to_signed(-141240030, 32), to_signed(-141444126, 32), to_signed(-141648217, 32), to_signed(-141852302, 32),
     to_signed(-142056382, 32), to_signed(-142260457, 32), to_signed(-142464527, 32), to_signed(-142668592, 32),
     to_signed(-142872651, 32), to_signed(-143076705, 32), to_signed(-143280754, 32), to_signed(-143484797, 32),
     to_signed(-143688835, 32), to_signed(-143892868, 32), to_signed(-144096896, 32), to_signed(-144300918, 32),
     to_signed(-144504935, 32), to_signed(-144708947, 32), to_signed(-144912954, 32), to_signed(-145116955, 32),
     to_signed(-145320950, 32), to_signed(-145524941, 32), to_signed(-145728926, 32), to_signed(-145932906, 32),
     to_signed(-146136880, 32), to_signed(-146340849, 32), to_signed(-146544812, 32), to_signed(-146748771, 32),
     to_signed(-146952723, 32), to_signed(-147156671, 32), to_signed(-147360613, 32), to_signed(-147564549, 32),
     to_signed(-147768480, 32), to_signed(-147972406, 32), to_signed(-148176326, 32), to_signed(-148380241, 32),
     to_signed(-148584150, 32), to_signed(-148788054, 32), to_signed(-148991953, 32), to_signed(-149195846, 32),
     to_signed(-149399733, 32), to_signed(-149603615, 32), to_signed(-149807492, 32), to_signed(-150011363, 32),
     to_signed(-150215228, 32), to_signed(-150419088, 32), to_signed(-150622942, 32), to_signed(-150826791, 32),
     to_signed(-151030634, 32), to_signed(-151234472, 32), to_signed(-151438304, 32), to_signed(-151642131, 32),
     to_signed(-151845952, 32), to_signed(-152049768, 32), to_signed(-152253577, 32), to_signed(-152457382, 32),
     to_signed(-152661180, 32), to_signed(-152864973, 32), to_signed(-153068761, 32), to_signed(-153272543, 32),
     to_signed(-153476319, 32), to_signed(-153680089, 32), to_signed(-153883854, 32), to_signed(-154087613, 32),
     to_signed(-154291367, 32), to_signed(-154495115, 32), to_signed(-154698857, 32), to_signed(-154902594, 32),
     to_signed(-155106324, 32), to_signed(-155310050, 32), to_signed(-155513769, 32), to_signed(-155717483, 32),
     to_signed(-155921191, 32), to_signed(-156124893, 32), to_signed(-156328589, 32), to_signed(-156532280, 32),
     to_signed(-156735965, 32), to_signed(-156939644, 32), to_signed(-157143318, 32), to_signed(-157346985, 32),
     to_signed(-157550647, 32), to_signed(-157754303, 32), to_signed(-157957954, 32), to_signed(-158161598, 32),
     to_signed(-158365237, 32), to_signed(-158568870, 32), to_signed(-158772497, 32), to_signed(-158976118, 32),
     to_signed(-159179733, 32), to_signed(-159383343, 32), to_signed(-159586946, 32), to_signed(-159790544, 32),
     to_signed(-159994136, 32), to_signed(-160197722, 32), to_signed(-160401302, 32), to_signed(-160604876, 32),
     to_signed(-160808445, 32), to_signed(-161012007, 32), to_signed(-161215564, 32), to_signed(-161419114, 32),
     to_signed(-161622659, 32), to_signed(-161826197, 32), to_signed(-162029730, 32), to_signed(-162233257, 32),
     to_signed(-162436778, 32), to_signed(-162640292, 32), to_signed(-162843801, 32), to_signed(-163047304, 32),
     to_signed(-163250801, 32), to_signed(-163454292, 32), to_signed(-163657777, 32), to_signed(-163861256, 32),
     to_signed(-164064728, 32), to_signed(-164268195, 32), to_signed(-164471656, 32), to_signed(-164675111, 32),
     to_signed(-164878559, 32), to_signed(-165082002, 32), to_signed(-165285438, 32), to_signed(-165488869, 32),
     to_signed(-165692293, 32), to_signed(-165895711, 32), to_signed(-166099124, 32), to_signed(-166302530, 32),
     to_signed(-166505929, 32), to_signed(-166709323, 32), to_signed(-166912711, 32), to_signed(-167116093, 32),
     to_signed(-167319468, 32), to_signed(-167522837, 32), to_signed(-167726200, 32), to_signed(-167929557, 32),
     to_signed(-168132908, 32), to_signed(-168336252, 32), to_signed(-168539591, 32), to_signed(-168742923, 32),
     to_signed(-168946249, 32), to_signed(-169149569, 32), to_signed(-169352882, 32), to_signed(-169556190, 32),
     to_signed(-169759491, 32), to_signed(-169962786, 32), to_signed(-170166074, 32), to_signed(-170369357, 32),
     to_signed(-170572633, 32), to_signed(-170775902, 32), to_signed(-170979166, 32), to_signed(-171182423, 32),
     to_signed(-171385674, 32), to_signed(-171588919, 32), to_signed(-171792157, 32), to_signed(-171995389, 32),
     to_signed(-172198615, 32), to_signed(-172401834, 32), to_signed(-172605047, 32), to_signed(-172808254, 32),
     to_signed(-173011454, 32), to_signed(-173214648, 32), to_signed(-173417836, 32), to_signed(-173621017, 32),
     to_signed(-173824192, 32), to_signed(-174027360, 32), to_signed(-174230522, 32), to_signed(-174433678, 32),
     to_signed(-174636827, 32), to_signed(-174839970, 32), to_signed(-175043106, 32), to_signed(-175246236, 32),
     to_signed(-175449360, 32), to_signed(-175652477, 32), to_signed(-175855587, 32), to_signed(-176058691, 32),
     to_signed(-176261789, 32), to_signed(-176464880, 32), to_signed(-176667965, 32), to_signed(-176871043, 32),
     to_signed(-177074115, 32), to_signed(-177277180, 32), to_signed(-177480239, 32), to_signed(-177683291, 32),
     to_signed(-177886336, 32), to_signed(-178089375, 32), to_signed(-178292408, 32), to_signed(-178495434, 32),
     to_signed(-178698453, 32), to_signed(-178901466, 32), to_signed(-179104472, 32), to_signed(-179307472, 32),
     to_signed(-179510465, 32), to_signed(-179713451, 32), to_signed(-179916431, 32), to_signed(-180119405, 32),
     to_signed(-180322371, 32), to_signed(-180525331, 32), to_signed(-180728284, 32), to_signed(-180931231, 32),
     to_signed(-181134171, 32), to_signed(-181337105, 32), to_signed(-181540031, 32), to_signed(-181742951, 32),
     to_signed(-181945865, 32), to_signed(-182148771, 32), to_signed(-182351671, 32), to_signed(-182554565, 32),
     to_signed(-182757451, 32), to_signed(-182960331, 32), to_signed(-183163204, 32), to_signed(-183366071, 32),
     to_signed(-183568930, 32), to_signed(-183771783, 32), to_signed(-183974629, 32), to_signed(-184177469, 32),
     to_signed(-184380301, 32), to_signed(-184583127, 32), to_signed(-184785946, 32), to_signed(-184988758, 32),
     to_signed(-185191564, 32), to_signed(-185394362, 32), to_signed(-185597154, 32), to_signed(-185799939, 32),
     to_signed(-186002717, 32), to_signed(-186205489, 32), to_signed(-186408253, 32), to_signed(-186611011, 32),
     to_signed(-186813762, 32), to_signed(-187016505, 32), to_signed(-187219242, 32), to_signed(-187421973, 32),
     to_signed(-187624696, 32), to_signed(-187827412, 32), to_signed(-188030122, 32), to_signed(-188232824, 32),
     to_signed(-188435520, 32), to_signed(-188638208, 32), to_signed(-188840890, 32), to_signed(-189043565, 32),
     to_signed(-189246233, 32), to_signed(-189448894, 32), to_signed(-189651548, 32), to_signed(-189854195, 32),
     to_signed(-190056834, 32), to_signed(-190259467, 32), to_signed(-190462093, 32), to_signed(-190664712, 32),
     to_signed(-190867324, 32), to_signed(-191069929, 32), to_signed(-191272527, 32), to_signed(-191475118, 32),
     to_signed(-191677702, 32), to_signed(-191880279, 32), to_signed(-192082849, 32), to_signed(-192285411, 32),
     to_signed(-192487967, 32), to_signed(-192690515, 32), to_signed(-192893057, 32), to_signed(-193095591, 32),
     to_signed(-193298119, 32), to_signed(-193500639, 32), to_signed(-193703152, 32), to_signed(-193905658, 32),
     to_signed(-194108156, 32), to_signed(-194310648, 32), to_signed(-194513133, 32), to_signed(-194715610, 32),
     to_signed(-194918080, 32), to_signed(-195120543, 32), to_signed(-195322999, 32), to_signed(-195525448, 32),
     to_signed(-195727889, 32), to_signed(-195930324, 32), to_signed(-196132751, 32), to_signed(-196335170, 32),
     to_signed(-196537583, 32), to_signed(-196739989, 32), to_signed(-196942387, 32), to_signed(-197144778, 32),
     to_signed(-197347161, 32), to_signed(-197549538, 32), to_signed(-197751907, 32), to_signed(-197954269, 32),
     to_signed(-198156624, 32), to_signed(-198358971, 32), to_signed(-198561311, 32), to_signed(-198763644, 32),
     to_signed(-198965969, 32), to_signed(-199168287, 32), to_signed(-199370598, 32), to_signed(-199572902, 32),
     to_signed(-199775198, 32), to_signed(-199977487, 32), to_signed(-200179768, 32), to_signed(-200382042, 32),
     to_signed(-200584309, 32), to_signed(-200786568, 32), to_signed(-200988820, 32), to_signed(-201191065, 32),
     to_signed(-201393302, 32), to_signed(-201595532, 32), to_signed(-201797754, 32), to_signed(-201999969, 32),
     to_signed(-202202177, 32), to_signed(-202404377, 32), to_signed(-202606569, 32), to_signed(-202808755, 32),
     to_signed(-203010932, 32), to_signed(-203213103, 32), to_signed(-203415265, 32), to_signed(-203617421, 32),
     to_signed(-203819569, 32), to_signed(-204021709, 32), to_signed(-204223842, 32), to_signed(-204425967, 32),
     to_signed(-204628085, 32), to_signed(-204830195, 32), to_signed(-205032298, 32), to_signed(-205234393, 32),
     to_signed(-205436481, 32), to_signed(-205638561, 32), to_signed(-205840633, 32), to_signed(-206042698, 32),
     to_signed(-206244756, 32), to_signed(-206446806, 32), to_signed(-206648848, 32), to_signed(-206850883, 32),
     to_signed(-207052910, 32), to_signed(-207254929, 32), to_signed(-207456941, 32), to_signed(-207658945, 32),
     to_signed(-207860942, 32), to_signed(-208062931, 32), to_signed(-208264912, 32), to_signed(-208466885, 32),
     to_signed(-208668851, 32), to_signed(-208870810, 32), to_signed(-209072760, 32), to_signed(-209274703, 32),
     to_signed(-209476638, 32), to_signed(-209678566, 32), to_signed(-209880485, 32), to_signed(-210082398, 32),
     to_signed(-210284302, 32), to_signed(-210486199, 32), to_signed(-210688087, 32), to_signed(-210889969, 32),
     to_signed(-211091842, 32), to_signed(-211293708, 32), to_signed(-211495565, 32), to_signed(-211697415, 32),
     to_signed(-211899258, 32), to_signed(-212101092, 32), to_signed(-212302919, 32), to_signed(-212504738, 32),
     to_signed(-212706549, 32), to_signed(-212908352, 32), to_signed(-213110148, 32), to_signed(-213311935, 32),
     to_signed(-213513715, 32), to_signed(-213715487, 32), to_signed(-213917251, 32), to_signed(-214119007, 32),
     to_signed(-214320755, 32), to_signed(-214522496, 32), to_signed(-214724228, 32), to_signed(-214925953, 32),
     to_signed(-215127670, 32), to_signed(-215329378, 32), to_signed(-215531079, 32), to_signed(-215732772, 32),
     to_signed(-215934457, 32), to_signed(-216136135, 32), to_signed(-216337804, 32), to_signed(-216539465, 32),
     to_signed(-216741118, 32), to_signed(-216942763, 32), to_signed(-217144401, 32), to_signed(-217346030, 32),
     to_signed(-217547651, 32), to_signed(-217749265, 32), to_signed(-217950870, 32), to_signed(-218152467, 32),
     to_signed(-218354057, 32), to_signed(-218555638, 32), to_signed(-218757211, 32), to_signed(-218958776, 32),
     to_signed(-219160334, 32), to_signed(-219361883, 32), to_signed(-219563424, 32), to_signed(-219764957, 32),
     to_signed(-219966481, 32), to_signed(-220167998, 32), to_signed(-220369507, 32), to_signed(-220571007, 32),
     to_signed(-220772500, 32), to_signed(-220973984, 32), to_signed(-221175461, 32), to_signed(-221376929, 32),
     to_signed(-221578389, 32), to_signed(-221779840, 32), to_signed(-221981284, 32), to_signed(-222182720, 32),
     to_signed(-222384147, 32), to_signed(-222585566, 32), to_signed(-222786977, 32), to_signed(-222988380, 32),
     to_signed(-223189774, 32), to_signed(-223391161, 32), to_signed(-223592539, 32), to_signed(-223793909, 32),
     to_signed(-223995270, 32), to_signed(-224196624, 32), to_signed(-224397969, 32), to_signed(-224599306, 32),
     to_signed(-224800635, 32), to_signed(-225001955, 32), to_signed(-225203267, 32), to_signed(-225404571, 32),
     to_signed(-225605867, 32), to_signed(-225807154, 32), to_signed(-226008433, 32), to_signed(-226209704, 32),
     to_signed(-226410966, 32), to_signed(-226612220, 32), to_signed(-226813466, 32), to_signed(-227014704, 32),
     to_signed(-227215933, 32), to_signed(-227417153, 32), to_signed(-227618366, 32), to_signed(-227819570, 32),
     to_signed(-228020765, 32), to_signed(-228221952, 32), to_signed(-228423131, 32), to_signed(-228624302, 32),
     to_signed(-228825464, 32), to_signed(-229026617, 32), to_signed(-229227762, 32), to_signed(-229428899, 32),
     to_signed(-229630027, 32), to_signed(-229831147, 32), to_signed(-230032259, 32), to_signed(-230233362, 32),
     to_signed(-230434456, 32), to_signed(-230635542, 32), to_signed(-230836620, 32), to_signed(-231037689, 32),
     to_signed(-231238749, 32), to_signed(-231439801, 32), to_signed(-231640845, 32), to_signed(-231841880, 32),
     to_signed(-232042906, 32), to_signed(-232243924, 32), to_signed(-232444934, 32), to_signed(-232645935, 32),
     to_signed(-232846927, 32), to_signed(-233047911, 32), to_signed(-233248886, 32), to_signed(-233449853, 32),
     to_signed(-233650811, 32), to_signed(-233851760, 32), to_signed(-234052701, 32), to_signed(-234253633, 32),
     to_signed(-234454557, 32), to_signed(-234655472, 32), to_signed(-234856378, 32), to_signed(-235057276, 32),
     to_signed(-235258165, 32), to_signed(-235459046, 32), to_signed(-235659918, 32), to_signed(-235860781, 32),
     to_signed(-236061635, 32), to_signed(-236262481, 32), to_signed(-236463318, 32), to_signed(-236664146, 32),
     to_signed(-236864966, 32), to_signed(-237065777, 32), to_signed(-237266579, 32), to_signed(-237467373, 32),
     to_signed(-237668158, 32), to_signed(-237868934, 32), to_signed(-238069701, 32), to_signed(-238270460, 32),
     to_signed(-238471210, 32), to_signed(-238671951, 32), to_signed(-238872683, 32), to_signed(-239073407, 32),
     to_signed(-239274121, 32), to_signed(-239474827, 32), to_signed(-239675524, 32), to_signed(-239876213, 32),
     to_signed(-240076892, 32), to_signed(-240277563, 32), to_signed(-240478225, 32), to_signed(-240678878, 32),
     to_signed(-240879522, 32), to_signed(-241080157, 32), to_signed(-241280783, 32), to_signed(-241481401, 32),
     to_signed(-241682010, 32), to_signed(-241882609, 32), to_signed(-242083200, 32), to_signed(-242283782, 32),
     to_signed(-242484355, 32), to_signed(-242684919, 32), to_signed(-242885475, 32), to_signed(-243086021, 32),
     to_signed(-243286558, 32), to_signed(-243487087, 32), to_signed(-243687606, 32), to_signed(-243888117, 32),
     to_signed(-244088618, 32), to_signed(-244289111, 32), to_signed(-244489594, 32), to_signed(-244690069, 32),
     to_signed(-244890535, 32), to_signed(-245090991, 32), to_signed(-245291439, 32), to_signed(-245491877, 32),
     to_signed(-245692307, 32), to_signed(-245892727, 32), to_signed(-246093139, 32), to_signed(-246293541, 32),
     to_signed(-246493935, 32), to_signed(-246694319, 32), to_signed(-246894694, 32), to_signed(-247095060, 32),
     to_signed(-247295417, 32), to_signed(-247495765, 32), to_signed(-247696104, 32), to_signed(-247896434, 32),
     to_signed(-248096755, 32), to_signed(-248297066, 32), to_signed(-248497369, 32), to_signed(-248697662, 32),
     to_signed(-248897946, 32), to_signed(-249098221, 32), to_signed(-249298487, 32), to_signed(-249498743, 32),
     to_signed(-249698991, 32), to_signed(-249899229, 32), to_signed(-250099458, 32), to_signed(-250299678, 32),
     to_signed(-250499889, 32), to_signed(-250700090, 32), to_signed(-250900283, 32), to_signed(-251100466, 32),
     to_signed(-251300640, 32), to_signed(-251500804, 32), to_signed(-251700959, 32), to_signed(-251901105, 32),
     to_signed(-252101242, 32), to_signed(-252301370, 32), to_signed(-252501488, 32), to_signed(-252701597, 32),
     to_signed(-252901697, 32), to_signed(-253101787, 32), to_signed(-253301868, 32), to_signed(-253501940, 32),
     to_signed(-253702003, 32), to_signed(-253902056, 32), to_signed(-254102099, 32), to_signed(-254302134, 32),
     to_signed(-254502159, 32), to_signed(-254702175, 32), to_signed(-254902181, 32), to_signed(-255102178, 32),
     to_signed(-255302166, 32), to_signed(-255502144, 32), to_signed(-255702113, 32), to_signed(-255902072, 32),
     to_signed(-256102022, 32), to_signed(-256301963, 32), to_signed(-256501894, 32), to_signed(-256701816, 32),
     to_signed(-256901728, 32), to_signed(-257101631, 32), to_signed(-257301525, 32), to_signed(-257501409, 32),
     to_signed(-257701283, 32), to_signed(-257901148, 32), to_signed(-258101004, 32), to_signed(-258300850, 32),
     to_signed(-258500686, 32), to_signed(-258700513, 32), to_signed(-258900331, 32), to_signed(-259100139, 32),
     to_signed(-259299937, 32), to_signed(-259499726, 32), to_signed(-259699506, 32), to_signed(-259899276, 32),
     to_signed(-260099036, 32), to_signed(-260298787, 32), to_signed(-260498528, 32), to_signed(-260698260, 32),
     to_signed(-260897982, 32), to_signed(-261097694, 32), to_signed(-261297397, 32), to_signed(-261497090, 32),
     to_signed(-261696774, 32), to_signed(-261896448, 32), to_signed(-262096112, 32), to_signed(-262295767, 32),
     to_signed(-262495412, 32), to_signed(-262695047, 32), to_signed(-262894673, 32), to_signed(-263094289, 32),
     to_signed(-263293896, 32), to_signed(-263493492, 32), to_signed(-263693079, 32), to_signed(-263892657, 32),
     to_signed(-264092224, 32), to_signed(-264291782, 32), to_signed(-264491331, 32), to_signed(-264690869, 32),
     to_signed(-264890398, 32), to_signed(-265089917, 32), to_signed(-265289426, 32), to_signed(-265488926, 32),
     to_signed(-265688415, 32), to_signed(-265887896, 32), to_signed(-266087366, 32), to_signed(-266286826, 32),
     to_signed(-266486277, 32), to_signed(-266685718, 32), to_signed(-266885149, 32), to_signed(-267084570, 32),
     to_signed(-267283981, 32), to_signed(-267483383, 32), to_signed(-267682775, 32), to_signed(-267882157, 32),
     to_signed(-268081529, 32), to_signed(-268280891, 32), to_signed(-268480243, 32), to_signed(-268679586, 32),
     to_signed(-268878918, 32), to_signed(-269078241, 32), to_signed(-269277554, 32), to_signed(-269476857, 32),
     to_signed(-269676150, 32), to_signed(-269875433, 32), to_signed(-270074706, 32), to_signed(-270273969, 32),
     to_signed(-270473223, 32), to_signed(-270672466, 32), to_signed(-270871700, 32), to_signed(-271070923, 32),
     to_signed(-271270136, 32), to_signed(-271469340, 32), to_signed(-271668533, 32), to_signed(-271867717, 32),
     to_signed(-272066891, 32), to_signed(-272266054, 32), to_signed(-272465208, 32), to_signed(-272664351, 32),
     to_signed(-272863485, 32), to_signed(-273062608, 32), to_signed(-273261722, 32), to_signed(-273460825, 32),
     to_signed(-273659918, 32), to_signed(-273859001, 32), to_signed(-274058075, 32), to_signed(-274257138, 32),
     to_signed(-274456191, 32), to_signed(-274655234, 32), to_signed(-274854267, 32), to_signed(-275053289, 32),
     to_signed(-275252302, 32), to_signed(-275451304, 32), to_signed(-275650297, 32), to_signed(-275849279, 32),
     to_signed(-276048251, 32), to_signed(-276247213, 32), to_signed(-276446165, 32), to_signed(-276645106, 32),
     to_signed(-276844038, 32), to_signed(-277042959, 32), to_signed(-277241870, 32), to_signed(-277440771, 32),
     to_signed(-277639662, 32), to_signed(-277838542, 32), to_signed(-278037413, 32), to_signed(-278236273, 32),
     to_signed(-278435122, 32), to_signed(-278633962, 32), to_signed(-278832791, 32), to_signed(-279031610, 32),
     to_signed(-279230419, 32), to_signed(-279429218, 32), to_signed(-279628006, 32), to_signed(-279826784, 32),
     to_signed(-280025552, 32), to_signed(-280224309, 32), to_signed(-280423056, 32), to_signed(-280621793, 32),
     to_signed(-280820520, 32), to_signed(-281019236, 32), to_signed(-281217942, 32), to_signed(-281416637, 32),
     to_signed(-281615322, 32), to_signed(-281813997, 32), to_signed(-282012662, 32), to_signed(-282211316, 32),
     to_signed(-282409959, 32), to_signed(-282608593, 32), to_signed(-282807215, 32), to_signed(-283005828, 32),
     to_signed(-283204430, 32), to_signed(-283403022, 32), to_signed(-283601603, 32), to_signed(-283800174, 32),
     to_signed(-283998734, 32), to_signed(-284197284, 32), to_signed(-284395824, 32), to_signed(-284594353, 32),
     to_signed(-284792871, 32), to_signed(-284991380, 32), to_signed(-285189877, 32), to_signed(-285388364, 32),
     to_signed(-285586841, 32), to_signed(-285785307, 32), to_signed(-285983763, 32), to_signed(-286182208, 32),
     to_signed(-286380643, 32), to_signed(-286579067, 32), to_signed(-286777480, 32), to_signed(-286975883, 32),
     to_signed(-287174276, 32), to_signed(-287372658, 32), to_signed(-287571029, 32), to_signed(-287769390, 32),
     to_signed(-287967740, 32), to_signed(-288166080, 32), to_signed(-288364409, 32), to_signed(-288562727, 32),
     to_signed(-288761035, 32), to_signed(-288959332, 32), to_signed(-289157619, 32), to_signed(-289355894, 32),
     to_signed(-289554160, 32), to_signed(-289752414, 32), to_signed(-289950658, 32), to_signed(-290148892, 32),
     to_signed(-290347114, 32), to_signed(-290545326, 32), to_signed(-290743528, 32), to_signed(-290941718, 32),
     to_signed(-291139898, 32), to_signed(-291338067, 32), to_signed(-291536226, 32), to_signed(-291734374, 32),
     to_signed(-291932511, 32), to_signed(-292130637, 32), to_signed(-292328753, 32), to_signed(-292526857, 32),
     to_signed(-292724951, 32), to_signed(-292923035, 32), to_signed(-293121107, 32), to_signed(-293319169, 32),
     to_signed(-293517220, 32), to_signed(-293715260, 32), to_signed(-293913290, 32), to_signed(-294111308, 32),
     to_signed(-294309316, 32), to_signed(-294507313, 32), to_signed(-294705299, 32), to_signed(-294903274, 32),
     to_signed(-295101239, 32), to_signed(-295299192, 32), to_signed(-295497135, 32), to_signed(-295695067, 32),
     to_signed(-295892988, 32), to_signed(-296090898, 32), to_signed(-296288797, 32), to_signed(-296486686, 32),
     to_signed(-296684563, 32), to_signed(-296882430, 32), to_signed(-297080285, 32), to_signed(-297278130, 32),
     to_signed(-297475964, 32), to_signed(-297673786, 32), to_signed(-297871598, 32), to_signed(-298069399, 32),
     to_signed(-298267189, 32), to_signed(-298464968, 32), to_signed(-298662736, 32), to_signed(-298860493, 32),
     to_signed(-299058239, 32), to_signed(-299255974, 32), to_signed(-299453698, 32), to_signed(-299651411, 32),
     to_signed(-299849113, 32), to_signed(-300046804, 32), to_signed(-300244484, 32), to_signed(-300442153, 32),
     to_signed(-300639811, 32), to_signed(-300837458, 32), to_signed(-301035094, 32), to_signed(-301232719, 32),
     to_signed(-301430332, 32), to_signed(-301627935, 32), to_signed(-301825526, 32), to_signed(-302023107, 32),
     to_signed(-302220676, 32), to_signed(-302418234, 32), to_signed(-302615781, 32), to_signed(-302813317, 32),
     to_signed(-303010842, 32), to_signed(-303208355, 32), to_signed(-303405858, 32), to_signed(-303603349, 32),
     to_signed(-303800829, 32), to_signed(-303998298, 32), to_signed(-304195756, 32), to_signed(-304393203, 32),
     to_signed(-304590638, 32), to_signed(-304788062, 32), to_signed(-304985475, 32), to_signed(-305182877, 32),
     to_signed(-305380268, 32), to_signed(-305577647, 32), to_signed(-305775015, 32), to_signed(-305972372, 32),
     to_signed(-306169718, 32), to_signed(-306367052, 32), to_signed(-306564375, 32), to_signed(-306761687, 32),
     to_signed(-306958988, 32), to_signed(-307156277, 32), to_signed(-307353555, 32), to_signed(-307550822, 32),
     to_signed(-307748077, 32), to_signed(-307945321, 32), to_signed(-308142554, 32), to_signed(-308339775, 32),
     to_signed(-308536985, 32), to_signed(-308734184, 32), to_signed(-308931371, 32), to_signed(-309128547, 32),
     to_signed(-309325712, 32), to_signed(-309522865, 32), to_signed(-309720007, 32), to_signed(-309917138, 32),
     to_signed(-310114257, 32), to_signed(-310311365, 32), to_signed(-310508461, 32), to_signed(-310705546, 32),
     to_signed(-310902619, 32), to_signed(-311099681, 32), to_signed(-311296732, 32), to_signed(-311493771, 32),
     to_signed(-311690799, 32), to_signed(-311887815, 32), to_signed(-312084820, 32), to_signed(-312281813, 32),
     to_signed(-312478795, 32), to_signed(-312675765, 32), to_signed(-312872724, 32), to_signed(-313069671, 32),
     to_signed(-313266607, 32), to_signed(-313463532, 32), to_signed(-313660444, 32), to_signed(-313857346, 32),
     to_signed(-314054235, 32), to_signed(-314251113, 32), to_signed(-314447980, 32), to_signed(-314644835, 32),
     to_signed(-314841679, 32), to_signed(-315038510, 32), to_signed(-315235331, 32), to_signed(-315432140, 32),
     to_signed(-315628937, 32), to_signed(-315825722, 32), to_signed(-316022496, 32), to_signed(-316219258, 32),
     to_signed(-316416009, 32), to_signed(-316612748, 32), to_signed(-316809475, 32), to_signed(-317006191, 32),
     to_signed(-317202895, 32), to_signed(-317399588, 32), to_signed(-317596268, 32), to_signed(-317792938, 32),
     to_signed(-317989595, 32), to_signed(-318186241, 32), to_signed(-318382875, 32), to_signed(-318579497, 32),
     to_signed(-318776108, 32), to_signed(-318972706, 32), to_signed(-319169293, 32), to_signed(-319365869, 32),
     to_signed(-319562433, 32), to_signed(-319758984, 32), to_signed(-319955525, 32), to_signed(-320152053, 32),
     to_signed(-320348570, 32), to_signed(-320545074, 32), to_signed(-320741568, 32), to_signed(-320938049, 32),
     to_signed(-321134518, 32), to_signed(-321330976, 32), to_signed(-321527422, 32), to_signed(-321723856, 32),
     to_signed(-321920278, 32), to_signed(-322116688, 32), to_signed(-322313087, 32), to_signed(-322509473, 32),
     to_signed(-322705848, 32), to_signed(-322902211, 32), to_signed(-323098562, 32), to_signed(-323294901, 32),
     to_signed(-323491229, 32), to_signed(-323687544, 32), to_signed(-323883848, 32), to_signed(-324080139, 32),
     to_signed(-324276419, 32), to_signed(-324472687, 32), to_signed(-324668942, 32), to_signed(-324865186, 32),
     to_signed(-325061418, 32), to_signed(-325257638, 32), to_signed(-325453846, 32), to_signed(-325650042, 32),
     to_signed(-325846226, 32), to_signed(-326042399, 32), to_signed(-326238559, 32), to_signed(-326434707, 32),
     to_signed(-326630843, 32), to_signed(-326826967, 32), to_signed(-327023079, 32), to_signed(-327219179, 32),
     to_signed(-327415267, 32), to_signed(-327611343, 32), to_signed(-327807407, 32), to_signed(-328003459, 32),
     to_signed(-328199499, 32), to_signed(-328395527, 32), to_signed(-328591543, 32), to_signed(-328787546, 32),
     to_signed(-328983538, 32), to_signed(-329179517, 32), to_signed(-329375485, 32), to_signed(-329571440, 32),
     to_signed(-329767383, 32), to_signed(-329963314, 32), to_signed(-330159233, 32), to_signed(-330355139, 32),
     to_signed(-330551034, 32), to_signed(-330746916, 32), to_signed(-330942787, 32), to_signed(-331138645, 32),
     to_signed(-331334491, 32), to_signed(-331530324, 32), to_signed(-331726146, 32), to_signed(-331921955, 32),
     to_signed(-332117752, 32), to_signed(-332313537, 32), to_signed(-332509310, 32), to_signed(-332705071, 32),
     to_signed(-332900819, 32), to_signed(-333096555, 32), to_signed(-333292279, 32), to_signed(-333487990, 32),
     to_signed(-333683689, 32), to_signed(-333879376, 32), to_signed(-334075051, 32), to_signed(-334270714, 32),
     to_signed(-334466364, 32), to_signed(-334662002, 32), to_signed(-334857627, 32), to_signed(-335053240, 32),
     to_signed(-335248841, 32), to_signed(-335444430, 32), to_signed(-335640006, 32), to_signed(-335835570, 32),
     to_signed(-336031121, 32), to_signed(-336226661, 32), to_signed(-336422188, 32), to_signed(-336617702, 32),
     to_signed(-336813204, 32), to_signed(-337008694, 32), to_signed(-337204171, 32), to_signed(-337399636, 32),
     to_signed(-337595089, 32), to_signed(-337790529, 32), to_signed(-337985956, 32), to_signed(-338181372, 32),
     to_signed(-338376774, 32), to_signed(-338572165, 32), to_signed(-338767543, 32), to_signed(-338962908, 32),
     to_signed(-339158261, 32), to_signed(-339353602, 32), to_signed(-339548930, 32), to_signed(-339744245, 32),
     to_signed(-339939549, 32), to_signed(-340134839, 32), to_signed(-340330117, 32), to_signed(-340525383, 32),
     to_signed(-340720636, 32), to_signed(-340915876, 32), to_signed(-341111104, 32), to_signed(-341306320, 32),
     to_signed(-341501523, 32), to_signed(-341696713, 32), to_signed(-341891891, 32), to_signed(-342087056, 32),
     to_signed(-342282209, 32), to_signed(-342477349, 32), to_signed(-342672476, 32), to_signed(-342867591, 32),
     to_signed(-343062693, 32), to_signed(-343257783, 32), to_signed(-343452860, 32), to_signed(-343647924, 32),
     to_signed(-343842976, 32), to_signed(-344038015, 32), to_signed(-344233042, 32), to_signed(-344428056, 32),
     to_signed(-344623057, 32), to_signed(-344818045, 32), to_signed(-345013021, 32), to_signed(-345207984, 32),
     to_signed(-345402934, 32), to_signed(-345597872, 32), to_signed(-345792797, 32), to_signed(-345987710, 32),
     to_signed(-346182609, 32), to_signed(-346377496, 32), to_signed(-346572370, 32), to_signed(-346767231, 32),
     to_signed(-346962080, 32), to_signed(-347156916, 32), to_signed(-347351739, 32), to_signed(-347546549, 32),
     to_signed(-347741347, 32), to_signed(-347936132, 32), to_signed(-348130904, 32), to_signed(-348325663, 32),
     to_signed(-348520409, 32), to_signed(-348715143, 32), to_signed(-348909863, 32), to_signed(-349104571, 32),
     to_signed(-349299266, 32), to_signed(-349493949, 32), to_signed(-349688618, 32), to_signed(-349883275, 32),
     to_signed(-350077918, 32), to_signed(-350272549, 32), to_signed(-350467167, 32), to_signed(-350661772, 32),
     to_signed(-350856364, 32), to_signed(-351050943, 32), to_signed(-351245510, 32), to_signed(-351440063, 32),
     to_signed(-351634604, 32), to_signed(-351829131, 32), to_signed(-352023646, 32), to_signed(-352218147, 32),
     to_signed(-352412636, 32), to_signed(-352607112, 32), to_signed(-352801575, 32), to_signed(-352996025, 32),
     to_signed(-353190461, 32), to_signed(-353384885, 32), to_signed(-353579296, 32), to_signed(-353773694, 32),
     to_signed(-353968079, 32), to_signed(-354162451, 32), to_signed(-354356810, 32), to_signed(-354551155, 32),
     to_signed(-354745488, 32), to_signed(-354939808, 32), to_signed(-355134115, 32), to_signed(-355328408, 32),
     to_signed(-355522689, 32), to_signed(-355716956, 32), to_signed(-355911211, 32), to_signed(-356105452, 32),
     to_signed(-356299680, 32), to_signed(-356493895, 32), to_signed(-356688097, 32), to_signed(-356882286, 32),
     to_signed(-357076462, 32), to_signed(-357270625, 32), to_signed(-357464774, 32), to_signed(-357658910, 32),
     to_signed(-357853034, 32), to_signed(-358047144, 32), to_signed(-358241241, 32), to_signed(-358435324, 32),
     to_signed(-358629395, 32), to_signed(-358823452, 32), to_signed(-359017496, 32), to_signed(-359211527, 32),
     to_signed(-359405545, 32), to_signed(-359599550, 32), to_signed(-359793541, 32), to_signed(-359987519, 32),
     to_signed(-360181484, 32), to_signed(-360375436, 32), to_signed(-360569374, 32), to_signed(-360763299, 32),
     to_signed(-360957211, 32), to_signed(-361151110, 32), to_signed(-361344995, 32), to_signed(-361538867, 32),
     to_signed(-361732726, 32), to_signed(-361926571, 32), to_signed(-362120403, 32), to_signed(-362314222, 32),
     to_signed(-362508027, 32), to_signed(-362701820, 32), to_signed(-362895598, 32), to_signed(-363089364, 32),
     to_signed(-363283116, 32), to_signed(-363476855, 32), to_signed(-363670580, 32), to_signed(-363864292, 32),
     to_signed(-364057991, 32), to_signed(-364251676, 32), to_signed(-364445348, 32), to_signed(-364639007, 32),
     to_signed(-364832652, 32), to_signed(-365026283, 32), to_signed(-365219902, 32), to_signed(-365413506, 32),
     to_signed(-365607098, 32), to_signed(-365800676, 32), to_signed(-365994240, 32), to_signed(-366187791, 32),
     to_signed(-366381329, 32), to_signed(-366574853, 32), to_signed(-366768363, 32), to_signed(-366961861, 32),
     to_signed(-367155344, 32), to_signed(-367348814, 32), to_signed(-367542271, 32), to_signed(-367735714, 32),
     to_signed(-367929144, 32), to_signed(-368122560, 32), to_signed(-368315962, 32), to_signed(-368509351, 32),
     to_signed(-368702727, 32), to_signed(-368896089, 32), to_signed(-369089437, 32), to_signed(-369282772, 32),
     to_signed(-369476093, 32), to_signed(-369669400, 32), to_signed(-369862694, 32), to_signed(-370055975, 32),
     to_signed(-370249242, 32), to_signed(-370442495, 32), to_signed(-370635734, 32), to_signed(-370828960, 32),
     to_signed(-371022173, 32), to_signed(-371215371, 32), to_signed(-371408556, 32), to_signed(-371601728, 32),
     to_signed(-371794885, 32), to_signed(-371988029, 32), to_signed(-372181160, 32), to_signed(-372374276, 32),
     to_signed(-372567379, 32), to_signed(-372760469, 32), to_signed(-372953544, 32), to_signed(-373146606, 32),
     to_signed(-373339654, 32), to_signed(-373532688, 32), to_signed(-373725709, 32), to_signed(-373918716, 32),
     to_signed(-374111709, 32), to_signed(-374304689, 32), to_signed(-374497654, 32), to_signed(-374690606, 32),
     to_signed(-374883544, 32), to_signed(-375076469, 32), to_signed(-375269379, 32), to_signed(-375462276, 32),
     to_signed(-375655159, 32), to_signed(-375848028, 32), to_signed(-376040883, 32), to_signed(-376233725, 32),
     to_signed(-376426553, 32), to_signed(-376619366, 32), to_signed(-376812166, 32), to_signed(-377004952, 32),
     to_signed(-377197725, 32), to_signed(-377390483, 32), to_signed(-377583228, 32), to_signed(-377775958, 32),
     to_signed(-377968675, 32), to_signed(-378161378, 32), to_signed(-378354067, 32), to_signed(-378546742, 32),
     to_signed(-378739403, 32), to_signed(-378932050, 32), to_signed(-379124683, 32), to_signed(-379317303, 32),
     to_signed(-379509908, 32), to_signed(-379702499, 32), to_signed(-379895077, 32), to_signed(-380087640, 32),
     to_signed(-380280190, 32), to_signed(-380472725, 32), to_signed(-380665247, 32), to_signed(-380857754, 32),
     to_signed(-381050248, 32), to_signed(-381242727, 32), to_signed(-381435193, 32), to_signed(-381627644, 32),
     to_signed(-381820082, 32), to_signed(-382012505, 32), to_signed(-382204915, 32), to_signed(-382397310, 32),
     to_signed(-382589691, 32), to_signed(-382782058, 32), to_signed(-382974412, 32), to_signed(-383166751, 32),
     to_signed(-383359076, 32), to_signed(-383551386, 32), to_signed(-383743683, 32), to_signed(-383935966, 32),
     to_signed(-384128234, 32), to_signed(-384320489, 32), to_signed(-384512729, 32), to_signed(-384704955, 32),
     to_signed(-384897167, 32), to_signed(-385089365, 32), to_signed(-385281549, 32), to_signed(-385473718, 32),
     to_signed(-385665873, 32), to_signed(-385858015, 32), to_signed(-386050142, 32), to_signed(-386242254, 32),
     to_signed(-386434353, 32), to_signed(-386626437, 32), to_signed(-386818508, 32), to_signed(-387010563, 32),
     to_signed(-387202605, 32), to_signed(-387394633, 32), to_signed(-387586646, 32), to_signed(-387778645, 32),
     to_signed(-387970630, 32), to_signed(-388162600, 32), to_signed(-388354556, 32), to_signed(-388546498, 32),
     to_signed(-388738426, 32), to_signed(-388930339, 32), to_signed(-389122238, 32), to_signed(-389314123, 32),
     to_signed(-389505993, 32), to_signed(-389697849, 32), to_signed(-389889691, 32), to_signed(-390081518, 32),
     to_signed(-390273331, 32), to_signed(-390465130, 32), to_signed(-390656915, 32), to_signed(-390848685, 32),
     to_signed(-391040440, 32), to_signed(-391232181, 32), to_signed(-391423908, 32), to_signed(-391615621, 32),
     to_signed(-391807319, 32), to_signed(-391999003, 32), to_signed(-392190672, 32), to_signed(-392382327, 32),
     to_signed(-392573967, 32), to_signed(-392765593, 32), to_signed(-392957205, 32), to_signed(-393148802, 32),
     to_signed(-393340384, 32), to_signed(-393531953, 32), to_signed(-393723506, 32), to_signed(-393915046, 32),
     to_signed(-394106570, 32), to_signed(-394298081, 32), to_signed(-394489576, 32), to_signed(-394681058, 32),
     to_signed(-394872524, 32), to_signed(-395063977, 32), to_signed(-395255414, 32), to_signed(-395446837, 32),
     to_signed(-395638246, 32), to_signed(-395829640, 32), to_signed(-396021020, 32), to_signed(-396212385, 32),
     to_signed(-396403735, 32), to_signed(-396595071, 32), to_signed(-396786392, 32), to_signed(-396977699, 32),
     to_signed(-397168991, 32), to_signed(-397360268, 32), to_signed(-397551531, 32), to_signed(-397742779, 32),
     to_signed(-397934013, 32), to_signed(-398125232, 32), to_signed(-398316436, 32), to_signed(-398507626, 32),
     to_signed(-398698801, 32), to_signed(-398889962, 32), to_signed(-399081107, 32), to_signed(-399272238, 32),
     to_signed(-399463355, 32), to_signed(-399654456, 32), to_signed(-399845543, 32), to_signed(-400036616, 32),
     to_signed(-400227673, 32), to_signed(-400418716, 32), to_signed(-400609744, 32), to_signed(-400800758, 32),
     to_signed(-400991756, 32), to_signed(-401182740, 32), to_signed(-401373709, 32), to_signed(-401564664, 32),
     to_signed(-401755603, 32), to_signed(-401946528, 32), to_signed(-402137438, 32), to_signed(-402328334, 32),
     to_signed(-402519214, 32), to_signed(-402710080, 32), to_signed(-402900931, 32), to_signed(-403091767, 32),
     to_signed(-403282588, 32), to_signed(-403473395, 32), to_signed(-403664186, 32), to_signed(-403854963, 32),
     to_signed(-404045725, 32), to_signed(-404236472, 32), to_signed(-404427204, 32), to_signed(-404617922, 32),
     to_signed(-404808624, 32), to_signed(-404999312, 32), to_signed(-405189985, 32), to_signed(-405380642, 32),
     to_signed(-405571285, 32), to_signed(-405761913, 32), to_signed(-405952526, 32), to_signed(-406143124, 32),
     to_signed(-406333708, 32), to_signed(-406524276, 32), to_signed(-406714829, 32), to_signed(-406905368, 32),
     to_signed(-407095891, 32), to_signed(-407286400, 32), to_signed(-407476893, 32), to_signed(-407667371, 32),
     to_signed(-407857835, 32), to_signed(-408048283, 32), to_signed(-408238717, 32), to_signed(-408429135, 32),
     to_signed(-408619539, 32), to_signed(-408809927, 32), to_signed(-409000301, 32), to_signed(-409190659, 32),
     to_signed(-409381002, 32), to_signed(-409571331, 32), to_signed(-409761644, 32), to_signed(-409951942, 32),
     to_signed(-410142225, 32), to_signed(-410332493, 32), to_signed(-410522746, 32), to_signed(-410712984, 32),
     to_signed(-410903207, 32), to_signed(-411093414, 32), to_signed(-411283607, 32), to_signed(-411473784, 32),
     to_signed(-411663946, 32), to_signed(-411854094, 32), to_signed(-412044226, 32), to_signed(-412234342, 32),
     to_signed(-412424444, 32), to_signed(-412614530, 32), to_signed(-412804602, 32), to_signed(-412994658, 32),
     to_signed(-413184699, 32), to_signed(-413374725, 32), to_signed(-413564735, 32), to_signed(-413754731, 32),
     to_signed(-413944711, 32), to_signed(-414134676, 32), to_signed(-414324625, 32), to_signed(-414514560, 32),
     to_signed(-414704479, 32), to_signed(-414894383, 32), to_signed(-415084272, 32), to_signed(-415274145, 32),
     to_signed(-415464004, 32), to_signed(-415653847, 32), to_signed(-415843674, 32), to_signed(-416033487, 32),
     to_signed(-416223284, 32), to_signed(-416413065, 32), to_signed(-416602832, 32), to_signed(-416792583, 32),
     to_signed(-416982319, 32), to_signed(-417172039, 32), to_signed(-417361744, 32), to_signed(-417551434, 32),
     to_signed(-417741109, 32), to_signed(-417930768, 32), to_signed(-418120411, 32), to_signed(-418310040, 32),
     to_signed(-418499653, 32), to_signed(-418689250, 32), to_signed(-418878833, 32), to_signed(-419068399, 32),
     to_signed(-419257951, 32), to_signed(-419447487, 32), to_signed(-419637007, 32), to_signed(-419826512, 32),
     to_signed(-420016002, 32), to_signed(-420205476, 32), to_signed(-420394935, 32), to_signed(-420584378, 32),
     to_signed(-420773806, 32), to_signed(-420963219, 32), to_signed(-421152615, 32), to_signed(-421341997, 32),
     to_signed(-421531363, 32), to_signed(-421720713, 32), to_signed(-421910048, 32), to_signed(-422099368, 32),
     to_signed(-422288671, 32), to_signed(-422477960, 32), to_signed(-422667233, 32), to_signed(-422856490, 32),
     to_signed(-423045732, 32), to_signed(-423234958, 32), to_signed(-423424169, 32), to_signed(-423613364, 32),
     to_signed(-423802543, 32), to_signed(-423991707, 32), to_signed(-424180855, 32), to_signed(-424369988, 32),
     to_signed(-424559105, 32), to_signed(-424748207, 32), to_signed(-424937293, 32), to_signed(-425126363, 32),
     to_signed(-425315418, 32), to_signed(-425504457, 32), to_signed(-425693480, 32), to_signed(-425882488, 32),
     to_signed(-426071480, 32), to_signed(-426260456, 32), to_signed(-426449417, 32), to_signed(-426638362, 32),
     to_signed(-426827291, 32), to_signed(-427016205, 32), to_signed(-427205103, 32), to_signed(-427393985, 32),
     to_signed(-427582852, 32), to_signed(-427771702, 32), to_signed(-427960537, 32), to_signed(-428149357, 32),
     to_signed(-428338160, 32), to_signed(-428526948, 32), to_signed(-428715720, 32), to_signed(-428904477, 32),
     to_signed(-429093217, 32), to_signed(-429281942, 32), to_signed(-429470651, 32), to_signed(-429659344, 32),
     to_signed(-429848022, 32), to_signed(-430036683, 32), to_signed(-430225329, 32), to_signed(-430413959, 32),
     to_signed(-430602573, 32), to_signed(-430791172, 32), to_signed(-430979754, 32), to_signed(-431168321, 32),
     to_signed(-431356872, 32), to_signed(-431545406, 32), to_signed(-431733926, 32), to_signed(-431922429, 32),
     to_signed(-432110916, 32), to_signed(-432299387, 32), to_signed(-432487843, 32), to_signed(-432676283, 32),
     to_signed(-432864706, 32), to_signed(-433053114, 32), to_signed(-433241506, 32), to_signed(-433429882, 32),
     to_signed(-433618242, 32), to_signed(-433806586, 32), to_signed(-433994914, 32), to_signed(-434183226, 32),
     to_signed(-434371523, 32), to_signed(-434559803, 32), to_signed(-434748067, 32), to_signed(-434936315, 32),
     to_signed(-435124548, 32), to_signed(-435312764, 32), to_signed(-435500964, 32), to_signed(-435689148, 32),
     to_signed(-435877317, 32), to_signed(-436065469, 32), to_signed(-436253605, 32), to_signed(-436441725, 32),
     to_signed(-436629829, 32), to_signed(-436817917, 32), to_signed(-437005989, 32), to_signed(-437194045, 32),
     to_signed(-437382085, 32), to_signed(-437570109, 32), to_signed(-437758117, 32), to_signed(-437946108, 32),
     to_signed(-438134084, 32), to_signed(-438322043, 32), to_signed(-438509986, 32), to_signed(-438697913, 32),
     to_signed(-438885824, 32), to_signed(-439073719, 32), to_signed(-439261598, 32), to_signed(-439449461, 32),
     to_signed(-439637307, 32), to_signed(-439825137, 32), to_signed(-440012951, 32), to_signed(-440200749, 32),
     to_signed(-440388531, 32), to_signed(-440576297, 32), to_signed(-440764046, 32), to_signed(-440951779, 32),
     to_signed(-441139496, 32), to_signed(-441327197, 32), to_signed(-441514881, 32), to_signed(-441702549, 32),
     to_signed(-441890201, 32), to_signed(-442077837, 32), to_signed(-442265456, 32), to_signed(-442453060, 32),
     to_signed(-442640647, 32), to_signed(-442828217, 32), to_signed(-443015772, 32), to_signed(-443203310, 32),
     to_signed(-443390832, 32), to_signed(-443578337, 32), to_signed(-443765826, 32), to_signed(-443953299, 32),
     to_signed(-444140756, 32), to_signed(-444328196, 32), to_signed(-444515620, 32), to_signed(-444703028, 32),
     to_signed(-444890419, 32), to_signed(-445077794, 32), to_signed(-445265152, 32), to_signed(-445452494, 32),
     to_signed(-445639820, 32), to_signed(-445827129, 32), to_signed(-446014422, 32), to_signed(-446201699, 32),
     to_signed(-446388959, 32), to_signed(-446576203, 32), to_signed(-446763430, 32), to_signed(-446950641, 32),
     to_signed(-447137835, 32), to_signed(-447325013, 32), to_signed(-447512175, 32), to_signed(-447699320, 32),
     to_signed(-447886449, 32), to_signed(-448073561, 32), to_signed(-448260657, 32), to_signed(-448447736, 32),
     to_signed(-448634799, 32), to_signed(-448821845, 32), to_signed(-449008875, 32), to_signed(-449195888, 32),
     to_signed(-449382885, 32), to_signed(-449569865, 32), to_signed(-449756829, 32), to_signed(-449943776, 32),
     to_signed(-450130706, 32), to_signed(-450317620, 32), to_signed(-450504518, 32), to_signed(-450691399, 32),
     to_signed(-450878263, 32), to_signed(-451065111, 32), to_signed(-451251942, 32), to_signed(-451438757, 32),
     to_signed(-451625555, 32), to_signed(-451812336, 32), to_signed(-451999101, 32), to_signed(-452185849, 32),
     to_signed(-452372581, 32), to_signed(-452559296, 32), to_signed(-452745994, 32), to_signed(-452932676, 32),
     to_signed(-453119340, 32), to_signed(-453305989, 32), to_signed(-453492620, 32), to_signed(-453679235, 32),
     to_signed(-453865834, 32), to_signed(-454052415, 32), to_signed(-454238980, 32), to_signed(-454425528, 32),
     to_signed(-454612060, 32), to_signed(-454798575, 32), to_signed(-454985073, 32), to_signed(-455171554, 32),
     to_signed(-455358019, 32), to_signed(-455544467, 32), to_signed(-455730898, 32), to_signed(-455917312, 32),
     to_signed(-456103710, 32), to_signed(-456290091, 32), to_signed(-456476455, 32), to_signed(-456662802, 32),
     to_signed(-456849132, 32), to_signed(-457035446, 32), to_signed(-457221743, 32), to_signed(-457408023, 32),
     to_signed(-457594286, 32), to_signed(-457780533, 32), to_signed(-457966762, 32), to_signed(-458152975, 32),
     to_signed(-458339171, 32), to_signed(-458525350, 32), to_signed(-458711512, 32), to_signed(-458897657, 32),
     to_signed(-459083786, 32), to_signed(-459269897, 32), to_signed(-459455992, 32), to_signed(-459642070, 32),
     to_signed(-459828131, 32), to_signed(-460014175, 32), to_signed(-460200202, 32), to_signed(-460386212, 32),
     to_signed(-460572205, 32), to_signed(-460758182, 32), to_signed(-460944141, 32), to_signed(-461130083, 32),
     to_signed(-461316009, 32), to_signed(-461501917, 32), to_signed(-461687809, 32), to_signed(-461873683, 32),
     to_signed(-462059541, 32), to_signed(-462245382, 32), to_signed(-462431205, 32), to_signed(-462617012, 32),
     to_signed(-462802801, 32), to_signed(-462988574, 32), to_signed(-463174329, 32), to_signed(-463360068, 32),
     to_signed(-463545789, 32), to_signed(-463731494, 32), to_signed(-463917181, 32), to_signed(-464102852, 32),
     to_signed(-464288505, 32), to_signed(-464474141, 32), to_signed(-464659760, 32), to_signed(-464845362, 32),
     to_signed(-465030947, 32), to_signed(-465216515, 32), to_signed(-465402066, 32), to_signed(-465587599, 32),
     to_signed(-465773116, 32), to_signed(-465958615, 32), to_signed(-466144097, 32), to_signed(-466329562, 32),
     to_signed(-466515010, 32), to_signed(-466700441, 32), to_signed(-466885855, 32), to_signed(-467071251, 32),
     to_signed(-467256631, 32), to_signed(-467441993, 32), to_signed(-467627338, 32), to_signed(-467812665, 32),
     to_signed(-467997976, 32), to_signed(-468183269, 32), to_signed(-468368545, 32), to_signed(-468553804, 32),
     to_signed(-468739046, 32), to_signed(-468924271, 32), to_signed(-469109478, 32), to_signed(-469294668, 32),
     to_signed(-469479840, 32), to_signed(-469664996, 32), to_signed(-469850134, 32), to_signed(-470035255, 32),
     to_signed(-470220358, 32), to_signed(-470405445, 32), to_signed(-470590514, 32), to_signed(-470775566, 32),
     to_signed(-470960600, 32), to_signed(-471145617, 32), to_signed(-471330617, 32), to_signed(-471515599, 32),
     to_signed(-471700564, 32), to_signed(-471885512, 32), to_signed(-472070443, 32), to_signed(-472255356, 32),
     to_signed(-472440251, 32), to_signed(-472625130, 32), to_signed(-472809991, 32), to_signed(-472994834, 32),
     to_signed(-473179660, 32), to_signed(-473364469, 32), to_signed(-473549261, 32), to_signed(-473734035, 32),
     to_signed(-473918791, 32), to_signed(-474103530, 32), to_signed(-474288252, 32), to_signed(-474472956, 32),
     to_signed(-474657643, 32), to_signed(-474842312, 32), to_signed(-475026964, 32), to_signed(-475211599, 32),
     to_signed(-475396216, 32), to_signed(-475580815, 32), to_signed(-475765397, 32), to_signed(-475949962, 32),
     to_signed(-476134509, 32), to_signed(-476319038, 32), to_signed(-476503550, 32), to_signed(-476688045, 32),
     to_signed(-476872522, 32), to_signed(-477056981, 32), to_signed(-477241423, 32), to_signed(-477425847, 32),
     to_signed(-477610254, 32), to_signed(-477794643, 32), to_signed(-477979015, 32), to_signed(-478163369, 32),
     to_signed(-478347705, 32), to_signed(-478532024, 32), to_signed(-478716326, 32), to_signed(-478900609, 32),
     to_signed(-479084875, 32), to_signed(-479269124, 32), to_signed(-479453355, 32), to_signed(-479637568, 32),
     to_signed(-479821764, 32), to_signed(-480005941, 32), to_signed(-480190102, 32), to_signed(-480374244, 32),
     to_signed(-480558369, 32), to_signed(-480742477, 32), to_signed(-480926566, 32), to_signed(-481110638, 32),
     to_signed(-481294693, 32), to_signed(-481478729, 32), to_signed(-481662748, 32), to_signed(-481846749, 32),
     to_signed(-482030733, 32), to_signed(-482214698, 32), to_signed(-482398646, 32), to_signed(-482582577, 32),
     to_signed(-482766489, 32), to_signed(-482950384, 32), to_signed(-483134261, 32), to_signed(-483318120, 32),
     to_signed(-483501962, 32), to_signed(-483685785, 32), to_signed(-483869591, 32), to_signed(-484053379, 32),
     to_signed(-484237150, 32), to_signed(-484420902, 32), to_signed(-484604637, 32), to_signed(-484788354, 32),
     to_signed(-484972053, 32), to_signed(-485155734, 32), to_signed(-485339398, 32), to_signed(-485523043, 32),
     to_signed(-485706671, 32), to_signed(-485890281, 32), to_signed(-486073873, 32), to_signed(-486257447, 32),
     to_signed(-486441003, 32), to_signed(-486624541, 32), to_signed(-486808062, 32), to_signed(-486991564, 32),
     to_signed(-487175049, 32), to_signed(-487358516, 32), to_signed(-487541965, 32), to_signed(-487725396, 32),
     to_signed(-487908809, 32), to_signed(-488092204, 32), to_signed(-488275581, 32), to_signed(-488458940, 32),
     to_signed(-488642281, 32), to_signed(-488825604, 32), to_signed(-489008909, 32), to_signed(-489192197, 32),
     to_signed(-489375466, 32), to_signed(-489558717, 32), to_signed(-489741950, 32), to_signed(-489925166, 32),
     to_signed(-490108363, 32), to_signed(-490291542, 32), to_signed(-490474703, 32), to_signed(-490657847, 32),
     to_signed(-490840972, 32), to_signed(-491024079, 32), to_signed(-491207168, 32), to_signed(-491390239, 32),
     to_signed(-491573292, 32), to_signed(-491756326, 32), to_signed(-491939343, 32), to_signed(-492122342, 32),
     to_signed(-492305322, 32), to_signed(-492488285, 32), to_signed(-492671229, 32), to_signed(-492854156, 32),
     to_signed(-493037064, 32), to_signed(-493219954, 32), to_signed(-493402826, 32), to_signed(-493585679, 32),
     to_signed(-493768515, 32), to_signed(-493951332, 32), to_signed(-494134132, 32), to_signed(-494316913, 32),
     to_signed(-494499676, 32), to_signed(-494682420, 32), to_signed(-494865147, 32), to_signed(-495047855, 32),
     to_signed(-495230545, 32), to_signed(-495413217, 32), to_signed(-495595871, 32), to_signed(-495778506, 32),
     to_signed(-495961124, 32), to_signed(-496143723, 32), to_signed(-496326304, 32), to_signed(-496508866, 32),
     to_signed(-496691410, 32), to_signed(-496873937, 32), to_signed(-497056444, 32), to_signed(-497238934, 32),
     to_signed(-497421405, 32), to_signed(-497603858, 32), to_signed(-497786293, 32), to_signed(-497968709, 32),
     to_signed(-498151107, 32), to_signed(-498333487, 32), to_signed(-498515848, 32), to_signed(-498698191, 32),
     to_signed(-498880516, 32), to_signed(-499062822, 32), to_signed(-499245110, 32), to_signed(-499427380, 32),
     to_signed(-499609631, 32), to_signed(-499791864, 32), to_signed(-499974079, 32), to_signed(-500156275, 32),
     to_signed(-500338453, 32), to_signed(-500520612, 32), to_signed(-500702753, 32), to_signed(-500884875, 32),
     to_signed(-501066980, 32), to_signed(-501249065, 32), to_signed(-501431133, 32), to_signed(-501613182, 32),
     to_signed(-501795212, 32), to_signed(-501977224, 32), to_signed(-502159217, 32), to_signed(-502341193, 32),
     to_signed(-502523149, 32), to_signed(-502705087, 32), to_signed(-502887007, 32), to_signed(-503068908, 32),
     to_signed(-503250791, 32), to_signed(-503432655, 32), to_signed(-503614500, 32), to_signed(-503796328, 32),
     to_signed(-503978136, 32), to_signed(-504159926, 32), to_signed(-504341698, 32), to_signed(-504523451, 32),
     to_signed(-504705185, 32), to_signed(-504886901, 32), to_signed(-505068598, 32), to_signed(-505250277, 32),
     to_signed(-505431937, 32), to_signed(-505613579, 32), to_signed(-505795202, 32), to_signed(-505976806, 32),
     to_signed(-506158392, 32), to_signed(-506339959, 32), to_signed(-506521508, 32), to_signed(-506703038, 32),
     to_signed(-506884549, 32), to_signed(-507066042, 32), to_signed(-507247516, 32), to_signed(-507428971, 32),
     to_signed(-507610408, 32), to_signed(-507791826, 32), to_signed(-507973225, 32), to_signed(-508154606, 32),
     to_signed(-508335968, 32), to_signed(-508517311, 32), to_signed(-508698636, 32), to_signed(-508879942, 32),
     to_signed(-509061229, 32), to_signed(-509242498, 32), to_signed(-509423748, 32), to_signed(-509604979, 32),
     to_signed(-509786191, 32), to_signed(-509967385, 32), to_signed(-510148559, 32), to_signed(-510329715, 32),
     to_signed(-510510853, 32), to_signed(-510691971, 32), to_signed(-510873071, 32), to_signed(-511054152, 32),
     to_signed(-511235214, 32), to_signed(-511416258, 32), to_signed(-511597282, 32), to_signed(-511778288, 32),
     to_signed(-511959275, 32), to_signed(-512140243, 32), to_signed(-512321192, 32), to_signed(-512502123, 32),
     to_signed(-512683035, 32), to_signed(-512863927, 32), to_signed(-513044801, 32), to_signed(-513225656, 32),
     to_signed(-513406493, 32), to_signed(-513587310, 32), to_signed(-513768108, 32), to_signed(-513948888, 32),
     to_signed(-514129648, 32), to_signed(-514310390, 32), to_signed(-514491113, 32), to_signed(-514671817, 32),
     to_signed(-514852502, 32), to_signed(-515033168, 32), to_signed(-515213815, 32), to_signed(-515394443, 32),
     to_signed(-515575053, 32), to_signed(-515755643, 32), to_signed(-515936214, 32), to_signed(-516116767, 32),
     to_signed(-516297300, 32), to_signed(-516477814, 32), to_signed(-516658310, 32), to_signed(-516838786, 32),
     to_signed(-517019243, 32), to_signed(-517199682, 32), to_signed(-517380101, 32), to_signed(-517560502, 32),
     to_signed(-517740883, 32), to_signed(-517921245, 32), to_signed(-518101588, 32), to_signed(-518281913, 32),
     to_signed(-518462218, 32), to_signed(-518642504, 32), to_signed(-518822771, 32), to_signed(-519003019, 32),
     to_signed(-519183248, 32), to_signed(-519363457, 32), to_signed(-519543648, 32), to_signed(-519723820, 32),
     to_signed(-519903972, 32), to_signed(-520084105, 32), to_signed(-520264220, 32), to_signed(-520444315, 32),
     to_signed(-520624391, 32), to_signed(-520804448, 32), to_signed(-520984485, 32), to_signed(-521164504, 32),
     to_signed(-521344503, 32), to_signed(-521524483, 32), to_signed(-521704444, 32), to_signed(-521884386, 32),
     to_signed(-522064309, 32), to_signed(-522244212, 32), to_signed(-522424096, 32), to_signed(-522603961, 32),
     to_signed(-522783807, 32), to_signed(-522963634, 32), to_signed(-523143441, 32), to_signed(-523323229, 32),
     to_signed(-523502998, 32), to_signed(-523682748, 32), to_signed(-523862478, 32), to_signed(-524042189, 32),
     to_signed(-524221881, 32), to_signed(-524401554, 32), to_signed(-524581207, 32), to_signed(-524760841, 32),
     to_signed(-524940456, 32), to_signed(-525120051, 32), to_signed(-525299627, 32), to_signed(-525479184, 32),
     to_signed(-525658722, 32), to_signed(-525838240, 32), to_signed(-526017739, 32), to_signed(-526197218, 32),
     to_signed(-526376678, 32), to_signed(-526556119, 32), to_signed(-526735541, 32), to_signed(-526914943, 32),
     to_signed(-527094325, 32), to_signed(-527273689, 32), to_signed(-527453033, 32), to_signed(-527632357, 32),
     to_signed(-527811662, 32), to_signed(-527990948, 32), to_signed(-528170214, 32), to_signed(-528349461, 32),
     to_signed(-528528689, 32), to_signed(-528707897, 32), to_signed(-528887085, 32), to_signed(-529066254, 32),
     to_signed(-529245404, 32), to_signed(-529424534, 32), to_signed(-529603645, 32), to_signed(-529782736, 32),
     to_signed(-529961808, 32), to_signed(-530140860, 32), to_signed(-530319893, 32), to_signed(-530498907, 32),
     to_signed(-530677900, 32), to_signed(-530856875, 32), to_signed(-531035830, 32), to_signed(-531214765, 32),
     to_signed(-531393681, 32), to_signed(-531572577, 32), to_signed(-531751453, 32), to_signed(-531930311, 32),
     to_signed(-532109148, 32), to_signed(-532287966, 32), to_signed(-532466765, 32), to_signed(-532645543, 32),
     to_signed(-532824303, 32), to_signed(-533003042, 32), to_signed(-533181762, 32), to_signed(-533360463, 32),
     to_signed(-533539144, 32), to_signed(-533717805, 32), to_signed(-533896447, 32), to_signed(-534075069, 32),
     to_signed(-534253671, 32), to_signed(-534432254, 32), to_signed(-534610817, 32), to_signed(-534789360, 32),
     to_signed(-534967884, 32), to_signed(-535146388, 32), to_signed(-535324872, 32), to_signed(-535503337, 32),
     to_signed(-535681782, 32), to_signed(-535860207, 32), to_signed(-536038613, 32), to_signed(-536216999, 32),
     to_signed(-536395365, 32), to_signed(-536573712, 32), to_signed(-536752038, 32), to_signed(-536930345, 32),
     to_signed(-537108633, 32), to_signed(-537286900, 32), to_signed(-537465148, 32), to_signed(-537643376, 32),
     to_signed(-537821584, 32), to_signed(-537999773, 32), to_signed(-538177942, 32), to_signed(-538356090, 32),
     to_signed(-538534220, 32), to_signed(-538712329, 32), to_signed(-538890418, 32), to_signed(-539068488, 32),
     to_signed(-539246538, 32), to_signed(-539424568, 32), to_signed(-539602578, 32), to_signed(-539780569, 32),
     to_signed(-539958539, 32), to_signed(-540136490, 32), to_signed(-540314421, 32), to_signed(-540492332, 32),
     to_signed(-540670223, 32), to_signed(-540848094, 32), to_signed(-541025945, 32), to_signed(-541203777, 32),
     to_signed(-541381588, 32), to_signed(-541559380, 32), to_signed(-541737151, 32), to_signed(-541914903, 32),
     to_signed(-542092635, 32), to_signed(-542270347, 32), to_signed(-542448039, 32), to_signed(-542625711, 32),
     to_signed(-542803363, 32), to_signed(-542980995, 32), to_signed(-543158607, 32), to_signed(-543336200, 32),
     to_signed(-543513772, 32), to_signed(-543691324, 32), to_signed(-543868856, 32), to_signed(-544046369, 32),
     to_signed(-544223861, 32), to_signed(-544401333, 32), to_signed(-544578785, 32), to_signed(-544756218, 32),
     to_signed(-544933630, 32), to_signed(-545111022, 32), to_signed(-545288394, 32), to_signed(-545465746, 32),
     to_signed(-545643078, 32), to_signed(-545820390, 32), to_signed(-545997682, 32), to_signed(-546174954, 32),
     to_signed(-546352205, 32), to_signed(-546529437, 32), to_signed(-546706649, 32), to_signed(-546883840, 32),
     to_signed(-547061011, 32), to_signed(-547238162, 32), to_signed(-547415294, 32), to_signed(-547592405, 32),
     to_signed(-547769495, 32), to_signed(-547946566, 32), to_signed(-548123617, 32), to_signed(-548300647, 32),
     to_signed(-548477657, 32), to_signed(-548654647, 32), to_signed(-548831617, 32), to_signed(-549008567, 32),
     to_signed(-549185496, 32), to_signed(-549362406, 32), to_signed(-549539295, 32), to_signed(-549716164, 32),
     to_signed(-549893013, 32), to_signed(-550069841, 32), to_signed(-550246649, 32), to_signed(-550423437, 32),
     to_signed(-550600205, 32), to_signed(-550776953, 32), to_signed(-550953680, 32), to_signed(-551130387, 32),
     to_signed(-551307074, 32), to_signed(-551483740, 32), to_signed(-551660387, 32), to_signed(-551837013, 32),
     to_signed(-552013618, 32), to_signed(-552190204, 32), to_signed(-552366769, 32), to_signed(-552543313, 32),
     to_signed(-552719838, 32), to_signed(-552896342, 32), to_signed(-553072826, 32), to_signed(-553249289, 32),
     to_signed(-553425732, 32), to_signed(-553602155, 32), to_signed(-553778558, 32), to_signed(-553954940, 32),
     to_signed(-554131301, 32), to_signed(-554307643, 32), to_signed(-554483964, 32), to_signed(-554660264, 32),
     to_signed(-554836544, 32), to_signed(-555012804, 32), to_signed(-555189044, 32), to_signed(-555365262, 32),
     to_signed(-555541461, 32), to_signed(-555717639, 32), to_signed(-555893797, 32), to_signed(-556069934, 32),
     to_signed(-556246051, 32), to_signed(-556422147, 32), to_signed(-556598223, 32), to_signed(-556774278, 32),
     to_signed(-556950313, 32), to_signed(-557126328, 32), to_signed(-557302322, 32), to_signed(-557478295, 32),
     to_signed(-557654248, 32), to_signed(-557830181, 32), to_signed(-558006093, 32), to_signed(-558181984, 32),
     to_signed(-558357855, 32), to_signed(-558533705, 32), to_signed(-558709535, 32), to_signed(-558885345, 32),
     to_signed(-559061133, 32), to_signed(-559236902, 32), to_signed(-559412649, 32), to_signed(-559588376, 32),
     to_signed(-559764083, 32), to_signed(-559939769, 32), to_signed(-560115434, 32), to_signed(-560291079, 32),
     to_signed(-560466703, 32), to_signed(-560642307, 32), to_signed(-560817890, 32), to_signed(-560993452, 32),
     to_signed(-561168994, 32), to_signed(-561344515, 32), to_signed(-561520015, 32), to_signed(-561695495, 32),
     to_signed(-561870954, 32), to_signed(-562046392, 32), to_signed(-562221810, 32), to_signed(-562397207, 32),
     to_signed(-562572584, 32), to_signed(-562747940, 32), to_signed(-562923275, 32), to_signed(-563098589, 32),
     to_signed(-563273883, 32), to_signed(-563449156, 32), to_signed(-563624408, 32), to_signed(-563799639, 32),
     to_signed(-563974850, 32), to_signed(-564150040, 32), to_signed(-564325210, 32), to_signed(-564500358, 32),
     to_signed(-564675486, 32), to_signed(-564850593, 32), to_signed(-565025679, 32), to_signed(-565200745, 32),
     to_signed(-565375790, 32), to_signed(-565550814, 32), to_signed(-565725817, 32), to_signed(-565900799, 32),
     to_signed(-566075761, 32), to_signed(-566250701, 32), to_signed(-566425621, 32), to_signed(-566600520, 32),
     to_signed(-566775399, 32), to_signed(-566950256, 32), to_signed(-567125093, 32), to_signed(-567299908, 32),
     to_signed(-567474703, 32), to_signed(-567649477, 32), to_signed(-567824230, 32), to_signed(-567998962, 32),
     to_signed(-568173674, 32), to_signed(-568348364, 32), to_signed(-568523034, 32), to_signed(-568697683, 32),
     to_signed(-568872310, 32), to_signed(-569046917, 32), to_signed(-569221503, 32), to_signed(-569396068, 32),
     to_signed(-569570612, 32), to_signed(-569745135, 32), to_signed(-569919637, 32), to_signed(-570094119, 32),
     to_signed(-570268579, 32), to_signed(-570443018, 32), to_signed(-570617437, 32), to_signed(-570791834, 32),
     to_signed(-570966210, 32), to_signed(-571140566, 32), to_signed(-571314900, 32), to_signed(-571489213, 32),
     to_signed(-571663506, 32), to_signed(-571837777, 32), to_signed(-572012027, 32), to_signed(-572186257, 32),
     to_signed(-572360465, 32), to_signed(-572534652, 32), to_signed(-572708818, 32), to_signed(-572882963, 32),
     to_signed(-573057087, 32), to_signed(-573231190, 32), to_signed(-573405272, 32), to_signed(-573579333, 32),
     to_signed(-573753372, 32), to_signed(-573927391, 32), to_signed(-574101389, 32), to_signed(-574275365, 32),
     to_signed(-574449320, 32), to_signed(-574623254, 32), to_signed(-574797167, 32), to_signed(-574971059, 32),
     to_signed(-575144930, 32), to_signed(-575318780, 32), to_signed(-575492608, 32), to_signed(-575666415, 32),
     to_signed(-575840202, 32), to_signed(-576013966, 32), to_signed(-576187710, 32), to_signed(-576361433, 32),
     to_signed(-576535134, 32), to_signed(-576708814, 32), to_signed(-576882473, 32), to_signed(-577056111, 32),
     to_signed(-577229728, 32), to_signed(-577403323, 32), to_signed(-577576897, 32), to_signed(-577750450, 32),
     to_signed(-577923982, 32), to_signed(-578097492, 32), to_signed(-578270981, 32), to_signed(-578444449, 32),
     to_signed(-578617896, 32), to_signed(-578791321, 32), to_signed(-578964725, 32), to_signed(-579138108, 32),
     to_signed(-579311470, 32), to_signed(-579484810, 32), to_signed(-579658129, 32), to_signed(-579831426, 32),
     to_signed(-580004702, 32), to_signed(-580177957, 32), to_signed(-580351191, 32), to_signed(-580524403, 32),
     to_signed(-580697594, 32), to_signed(-580870764, 32), to_signed(-581043912, 32), to_signed(-581217039, 32),
     to_signed(-581390144, 32), to_signed(-581563228, 32), to_signed(-581736291, 32), to_signed(-581909332, 32),
     to_signed(-582082352, 32), to_signed(-582255351, 32), to_signed(-582428328, 32), to_signed(-582601283, 32),
     to_signed(-582774218, 32), to_signed(-582947131, 32), to_signed(-583120022, 32), to_signed(-583292892, 32),
     to_signed(-583465740, 32), to_signed(-583638568, 32), to_signed(-583811373, 32), to_signed(-583984157, 32),
     to_signed(-584156920, 32), to_signed(-584329661, 32), to_signed(-584502381, 32), to_signed(-584675079, 32),
     to_signed(-584847756, 32), to_signed(-585020411, 32), to_signed(-585193045, 32), to_signed(-585365657, 32),
     to_signed(-585538248, 32), to_signed(-585710817, 32), to_signed(-585883365, 32), to_signed(-586055891, 32),
     to_signed(-586228395, 32), to_signed(-586400878, 32), to_signed(-586573340, 32), to_signed(-586745779, 32),
     to_signed(-586918198, 32), to_signed(-587090594, 32), to_signed(-587262969, 32), to_signed(-587435323, 32),
     to_signed(-587607655, 32), to_signed(-587779965, 32), to_signed(-587952254, 32), to_signed(-588124521, 32),
     to_signed(-588296766, 32), to_signed(-588468990, 32), to_signed(-588641192, 32), to_signed(-588813373, 32),
     to_signed(-588985532, 32), to_signed(-589157669, 32), to_signed(-589329785, 32), to_signed(-589501879, 32),
     to_signed(-589673951, 32), to_signed(-589846002, 32), to_signed(-590018030, 32), to_signed(-590190038, 32),
     to_signed(-590362023, 32), to_signed(-590533987, 32), to_signed(-590705929, 32), to_signed(-590877849, 32),
     to_signed(-591049748, 32), to_signed(-591221625, 32), to_signed(-591393480, 32), to_signed(-591565313, 32),
     to_signed(-591737125, 32), to_signed(-591908915, 32), to_signed(-592080683, 32), to_signed(-592252429, 32),
     to_signed(-592424154, 32), to_signed(-592595857, 32), to_signed(-592767538, 32), to_signed(-592939197, 32),
     to_signed(-593110835, 32), to_signed(-593282450, 32), to_signed(-593454044, 32), to_signed(-593625616, 32),
     to_signed(-593797166, 32), to_signed(-593968694, 32), to_signed(-594140201, 32), to_signed(-594311686, 32),
     to_signed(-594483148, 32), to_signed(-594654589, 32), to_signed(-594826008, 32), to_signed(-594997406, 32),
     to_signed(-595168781, 32), to_signed(-595340134, 32), to_signed(-595511466, 32), to_signed(-595682776, 32),
     to_signed(-595854063, 32), to_signed(-596025329, 32), to_signed(-596196573, 32), to_signed(-596367795, 32),
     to_signed(-596538995, 32), to_signed(-596710174, 32), to_signed(-596881330, 32), to_signed(-597052464, 32),
     to_signed(-597223576, 32), to_signed(-597394667, 32), to_signed(-597565735, 32), to_signed(-597736782, 32),
     to_signed(-597907806, 32), to_signed(-598078808, 32), to_signed(-598249789, 32), to_signed(-598420747, 32),
     to_signed(-598591684, 32), to_signed(-598762598, 32), to_signed(-598933491, 32), to_signed(-599104361, 32),
     to_signed(-599275210, 32), to_signed(-599446036, 32), to_signed(-599616840, 32), to_signed(-599787623, 32),
     to_signed(-599958383, 32), to_signed(-600129121, 32), to_signed(-600299837, 32), to_signed(-600470531, 32),
     to_signed(-600641203, 32), to_signed(-600811853, 32), to_signed(-600982481, 32), to_signed(-601153087, 32),
     to_signed(-601323670, 32), to_signed(-601494232, 32), to_signed(-601664771, 32), to_signed(-601835288, 32),
     to_signed(-602005783, 32), to_signed(-602176256, 32), to_signed(-602346707, 32), to_signed(-602517136, 32),
     to_signed(-602687543, 32), to_signed(-602857927, 32), to_signed(-603028289, 32), to_signed(-603198629, 32),
     to_signed(-603368947, 32), to_signed(-603539243, 32), to_signed(-603709516, 32), to_signed(-603879768, 32),
     to_signed(-604049997, 32), to_signed(-604220204, 32), to_signed(-604390388, 32), to_signed(-604560551, 32),
     to_signed(-604730691, 32), to_signed(-604900809, 32), to_signed(-605070905, 32), to_signed(-605240978, 32),
     to_signed(-605411029, 32), to_signed(-605581058, 32), to_signed(-605751065, 32), to_signed(-605921050, 32),
     to_signed(-606091012, 32), to_signed(-606260952, 32), to_signed(-606430869, 32), to_signed(-606600765, 32),
     to_signed(-606770638, 32), to_signed(-606940488, 32), to_signed(-607110317, 32), to_signed(-607280123, 32),
     to_signed(-607449906, 32), to_signed(-607619668, 32), to_signed(-607789407, 32), to_signed(-607959124, 32),
     to_signed(-608128818, 32), to_signed(-608298490, 32), to_signed(-608468140, 32), to_signed(-608637767, 32),
     to_signed(-608807372, 32), to_signed(-608976954, 32), to_signed(-609146514, 32), to_signed(-609316052, 32),
     to_signed(-609485567, 32), to_signed(-609655060, 32), to_signed(-609824531, 32), to_signed(-609993979, 32),
     to_signed(-610163404, 32), to_signed(-610332808, 32), to_signed(-610502188, 32), to_signed(-610671547, 32),
     to_signed(-610840882, 32), to_signed(-611010196, 32), to_signed(-611179487, 32), to_signed(-611348755, 32),
     to_signed(-611518001, 32), to_signed(-611687225, 32), to_signed(-611856426, 32), to_signed(-612025604, 32),
     to_signed(-612194760, 32), to_signed(-612363894, 32), to_signed(-612533005, 32), to_signed(-612702093, 32),
     to_signed(-612871159, 32), to_signed(-613040203, 32), to_signed(-613209223, 32), to_signed(-613378222, 32),
     to_signed(-613547198, 32), to_signed(-613716151, 32), to_signed(-613885081, 32), to_signed(-614053989, 32),
     to_signed(-614222875, 32), to_signed(-614391738, 32), to_signed(-614560578, 32), to_signed(-614729396, 32),
     to_signed(-614898191, 32), to_signed(-615066964, 32), to_signed(-615235714, 32), to_signed(-615404441, 32),
     to_signed(-615573145, 32), to_signed(-615741827, 32), to_signed(-615910487, 32), to_signed(-616079124, 32),
     to_signed(-616247738, 32), to_signed(-616416329, 32), to_signed(-616584898, 32), to_signed(-616753444, 32),
     to_signed(-616921967, 32), to_signed(-617090468, 32), to_signed(-617258946, 32), to_signed(-617427402, 32),
     to_signed(-617595834, 32), to_signed(-617764244, 32), to_signed(-617932631, 32), to_signed(-618100996, 32),
     to_signed(-618269338, 32), to_signed(-618437657, 32), to_signed(-618605953, 32), to_signed(-618774227, 32),
     to_signed(-618942478, 32), to_signed(-619110706, 32), to_signed(-619278911, 32), to_signed(-619447093, 32),
     to_signed(-619615253, 32), to_signed(-619783390, 32), to_signed(-619951504, 32), to_signed(-620119596, 32),
     to_signed(-620287664, 32), to_signed(-620455710, 32), to_signed(-620623733, 32), to_signed(-620791733, 32),
     to_signed(-620959711, 32), to_signed(-621127665, 32), to_signed(-621295597, 32), to_signed(-621463506, 32),
     to_signed(-621631392, 32), to_signed(-621799255, 32), to_signed(-621967095, 32), to_signed(-622134912, 32),
     to_signed(-622302707, 32), to_signed(-622470478, 32), to_signed(-622638227, 32), to_signed(-622805953, 32),
     to_signed(-622973656, 32), to_signed(-623141336, 32), to_signed(-623308993, 32), to_signed(-623476627, 32),
     to_signed(-623644239, 32), to_signed(-623811827, 32), to_signed(-623979393, 32), to_signed(-624146935, 32),
     to_signed(-624314455, 32), to_signed(-624481951, 32), to_signed(-624649425, 32), to_signed(-624816875, 32),
     to_signed(-624984303, 32), to_signed(-625151708, 32), to_signed(-625319090, 32), to_signed(-625486448, 32),
     to_signed(-625653784, 32), to_signed(-625821097, 32), to_signed(-625988387, 32), to_signed(-626155653, 32),
     to_signed(-626322897, 32), to_signed(-626490118, 32), to_signed(-626657315, 32), to_signed(-626824490, 32),
     to_signed(-626991641, 32), to_signed(-627158770, 32), to_signed(-627325875, 32), to_signed(-627492958, 32),
     to_signed(-627660017, 32), to_signed(-627827053, 32), to_signed(-627994066, 32), to_signed(-628161056, 32),
     to_signed(-628328023, 32), to_signed(-628494967, 32), to_signed(-628661888, 32), to_signed(-628828785, 32),
     to_signed(-628995660, 32), to_signed(-629162511, 32), to_signed(-629329340, 32), to_signed(-629496145, 32),
     to_signed(-629662927, 32), to_signed(-629829685, 32), to_signed(-629996421, 32), to_signed(-630163134, 32),
     to_signed(-630329823, 32), to_signed(-630496489, 32), to_signed(-630663132, 32), to_signed(-630829752, 32),
     to_signed(-630996348, 32), to_signed(-631162922, 32), to_signed(-631329472, 32), to_signed(-631495999, 32),
     to_signed(-631662503, 32), to_signed(-631828983, 32), to_signed(-631995440, 32), to_signed(-632161874, 32),
     to_signed(-632328285, 32), to_signed(-632494673, 32), to_signed(-632661037, 32), to_signed(-632827378, 32),
     to_signed(-632993696, 32), to_signed(-633159990, 32), to_signed(-633326262, 32), to_signed(-633492510, 32),
     to_signed(-633658734, 32), to_signed(-633824936, 32), to_signed(-633991114, 32), to_signed(-634157268, 32),
     to_signed(-634323400, 32), to_signed(-634489508, 32), to_signed(-634655593, 32), to_signed(-634821654, 32),
     to_signed(-634987692, 32), to_signed(-635153707, 32), to_signed(-635319698, 32), to_signed(-635485666, 32),
     to_signed(-635651611, 32), to_signed(-635817532, 32), to_signed(-635983430, 32), to_signed(-636149305, 32),
     to_signed(-636315156, 32), to_signed(-636480984, 32), to_signed(-636646788, 32), to_signed(-636812569, 32),
     to_signed(-636978327, 32), to_signed(-637144061, 32), to_signed(-637309771, 32), to_signed(-637475459, 32),
     to_signed(-637641122, 32), to_signed(-637806763, 32), to_signed(-637972380, 32), to_signed(-638137973, 32),
     to_signed(-638303543, 32), to_signed(-638469090, 32), to_signed(-638634613, 32), to_signed(-638800112, 32),
     to_signed(-638965588, 32), to_signed(-639131041, 32), to_signed(-639296470, 32), to_signed(-639461876, 32),
     to_signed(-639627258, 32), to_signed(-639792616, 32), to_signed(-639957951, 32), to_signed(-640123263, 32),
     to_signed(-640288551, 32), to_signed(-640453815, 32), to_signed(-640619056, 32), to_signed(-640784274, 32),
     to_signed(-640949467, 32), to_signed(-641114637, 32), to_signed(-641279784, 32), to_signed(-641444907, 32),
     to_signed(-641610007, 32), to_signed(-641775083, 32), to_signed(-641940135, 32), to_signed(-642105163, 32),
     to_signed(-642270169, 32), to_signed(-642435150, 32), to_signed(-642600108, 32), to_signed(-642765042, 32),
     to_signed(-642929953, 32), to_signed(-643094840, 32), to_signed(-643259703, 32), to_signed(-643424543, 32),
     to_signed(-643589359, 32), to_signed(-643754151, 32), to_signed(-643918920, 32), to_signed(-644083665, 32),
     to_signed(-644248386, 32), to_signed(-644413083, 32), to_signed(-644577757, 32), to_signed(-644742408, 32),
     to_signed(-644907034, 32), to_signed(-645071637, 32), to_signed(-645236216, 32), to_signed(-645400771, 32),
     to_signed(-645565303, 32), to_signed(-645729811, 32), to_signed(-645894295, 32), to_signed(-646058755, 32),
     to_signed(-646223192, 32), to_signed(-646387605, 32), to_signed(-646551994, 32), to_signed(-646716360, 32),
     to_signed(-646880701, 32), to_signed(-647045019, 32), to_signed(-647209313, 32), to_signed(-647373583, 32),
     to_signed(-647537830, 32), to_signed(-647702052, 32), to_signed(-647866251, 32), to_signed(-648030426, 32),
     to_signed(-648194577, 32), to_signed(-648358704, 32), to_signed(-648522808, 32), to_signed(-648686887, 32),
     to_signed(-648850943, 32), to_signed(-649014975, 32), to_signed(-649178983, 32), to_signed(-649342967, 32),
     to_signed(-649506928, 32), to_signed(-649670864, 32), to_signed(-649834777, 32), to_signed(-649998665, 32),
     to_signed(-650162530, 32), to_signed(-650326371, 32), to_signed(-650490188, 32), to_signed(-650653981, 32),
     to_signed(-650817750, 32), to_signed(-650981495, 32), to_signed(-651145216, 32), to_signed(-651308914, 32),
     to_signed(-651472587, 32), to_signed(-651636236, 32), to_signed(-651799862, 32), to_signed(-651963463, 32),
     to_signed(-652127041, 32), to_signed(-652290594, 32), to_signed(-652454124, 32), to_signed(-652617629, 32),
     to_signed(-652781111, 32), to_signed(-652944569, 32), to_signed(-653108002, 32), to_signed(-653271412, 32),
     to_signed(-653434797, 32), to_signed(-653598159, 32), to_signed(-653761496, 32), to_signed(-653924810, 32),
     to_signed(-654088099, 32), to_signed(-654251364, 32), to_signed(-654414606, 32), to_signed(-654577823, 32),
     to_signed(-654741016, 32), to_signed(-654904185, 32), to_signed(-655067330, 32), to_signed(-655230451, 32),
     to_signed(-655393548, 32), to_signed(-655556620, 32), to_signed(-655719669, 32), to_signed(-655882694, 32),
     to_signed(-656045694, 32), to_signed(-656208670, 32), to_signed(-656371622, 32), to_signed(-656534550, 32),
     to_signed(-656697454, 32), to_signed(-656860334, 32), to_signed(-657023190, 32), to_signed(-657186021, 32),
     to_signed(-657348828, 32), to_signed(-657511611, 32), to_signed(-657674370, 32), to_signed(-657837105, 32),
     to_signed(-657999816, 32), to_signed(-658162502, 32), to_signed(-658325164, 32), to_signed(-658487802, 32),
     to_signed(-658650416, 32), to_signed(-658813005, 32), to_signed(-658975571, 32), to_signed(-659138112, 32),
     to_signed(-659300629, 32), to_signed(-659463121, 32), to_signed(-659625590, 32), to_signed(-659788034, 32),
     to_signed(-659950454, 32), to_signed(-660112849, 32), to_signed(-660275220, 32), to_signed(-660437568, 32),
     to_signed(-660599890, 32), to_signed(-660762189, 32), to_signed(-660924463, 32), to_signed(-661086713, 32),
     to_signed(-661248938, 32), to_signed(-661411140, 32), to_signed(-661573317, 32), to_signed(-661735469, 32),
     to_signed(-661897597, 32), to_signed(-662059701, 32), to_signed(-662221781, 32), to_signed(-662383836, 32),
     to_signed(-662545867, 32), to_signed(-662707874, 32), to_signed(-662869856, 32), to_signed(-663031814, 32),
     to_signed(-663193747, 32), to_signed(-663355656, 32), to_signed(-663517541, 32), to_signed(-663679401, 32),
     to_signed(-663841237, 32), to_signed(-664003048, 32), to_signed(-664164835, 32), to_signed(-664326598, 32),
     to_signed(-664488336, 32), to_signed(-664650050, 32), to_signed(-664811739, 32), to_signed(-664973404, 32),
     to_signed(-665135044, 32), to_signed(-665296660, 32), to_signed(-665458252, 32), to_signed(-665619819, 32),
     to_signed(-665781362, 32), to_signed(-665942880, 32), to_signed(-666104373, 32), to_signed(-666265842, 32),
     to_signed(-666427287, 32), to_signed(-666588707, 32), to_signed(-666750103, 32), to_signed(-666911474, 32),
     to_signed(-667072820, 32), to_signed(-667234142, 32), to_signed(-667395440, 32), to_signed(-667556713, 32),
     to_signed(-667717961, 32), to_signed(-667879185, 32), to_signed(-668040385, 32), to_signed(-668201559, 32),
     to_signed(-668362709, 32), to_signed(-668523835, 32), to_signed(-668684936, 32), to_signed(-668846013, 32),
     to_signed(-669007064, 32), to_signed(-669168092, 32), to_signed(-669329094, 32), to_signed(-669490072, 32),
     to_signed(-669651026, 32), to_signed(-669811955, 32), to_signed(-669972859, 32), to_signed(-670133738, 32),
     to_signed(-670294593, 32), to_signed(-670455424, 32), to_signed(-670616229, 32), to_signed(-670777010, 32),
     to_signed(-670937767, 32), to_signed(-671098498, 32), to_signed(-671259205, 32), to_signed(-671419887, 32),
     to_signed(-671580545, 32), to_signed(-671741178, 32), to_signed(-671901786, 32), to_signed(-672062370, 32),
     to_signed(-672222928, 32), to_signed(-672383462, 32), to_signed(-672543972, 32), to_signed(-672704456, 32),
     to_signed(-672864916, 32), to_signed(-673025352, 32), to_signed(-673185762, 32), to_signed(-673346148, 32),
     to_signed(-673506508, 32), to_signed(-673666845, 32), to_signed(-673827156, 32), to_signed(-673987443, 32),
     to_signed(-674147704, 32), to_signed(-674307941, 32), to_signed(-674468154, 32), to_signed(-674628341, 32),
     to_signed(-674788504, 32), to_signed(-674948642, 32), to_signed(-675108755, 32), to_signed(-675268843, 32),
     to_signed(-675428906, 32), to_signed(-675588945, 32), to_signed(-675748958, 32), to_signed(-675908947, 32),
     to_signed(-676068911, 32), to_signed(-676228850, 32), to_signed(-676388765, 32), to_signed(-676548654, 32),
     to_signed(-676708518, 32), to_signed(-676868358, 32), to_signed(-677028173, 32), to_signed(-677187963, 32),
     to_signed(-677347728, 32), to_signed(-677507468, 32), to_signed(-677667183, 32), to_signed(-677826873, 32),
     to_signed(-677986538, 32), to_signed(-678146179, 32), to_signed(-678305794, 32), to_signed(-678465385, 32),
     to_signed(-678624950, 32), to_signed(-678784491, 32), to_signed(-678944007, 32), to_signed(-679103497, 32),
     to_signed(-679262963, 32), to_signed(-679422404, 32), to_signed(-679581820, 32), to_signed(-679741210, 32),
     to_signed(-679900576, 32), to_signed(-680059917, 32), to_signed(-680219233, 32), to_signed(-680378524, 32),
     to_signed(-680537789, 32), to_signed(-680697030, 32), to_signed(-680856246, 32), to_signed(-681015436, 32),
     to_signed(-681174602, 32), to_signed(-681333743, 32), to_signed(-681492858, 32), to_signed(-681651949, 32),
     to_signed(-681811014, 32), to_signed(-681970055, 32), to_signed(-682129070, 32), to_signed(-682288060, 32),
     to_signed(-682447025, 32), to_signed(-682605965, 32), to_signed(-682764880, 32), to_signed(-682923770, 32),
     to_signed(-683082635, 32), to_signed(-683241474, 32), to_signed(-683400289, 32), to_signed(-683559078, 32),
     to_signed(-683717842, 32), to_signed(-683876581, 32), to_signed(-684035295, 32), to_signed(-684193984, 32),
     to_signed(-684352648, 32), to_signed(-684511286, 32), to_signed(-684669900, 32), to_signed(-684828488, 32),
     to_signed(-684987051, 32), to_signed(-685145588, 32), to_signed(-685304101, 32), to_signed(-685462588, 32),
     to_signed(-685621051, 32), to_signed(-685779488, 32), to_signed(-685937899, 32), to_signed(-686096286, 32),
     to_signed(-686254647, 32), to_signed(-686412983, 32), to_signed(-686571294, 32), to_signed(-686729580, 32),
     to_signed(-686887840, 32), to_signed(-687046075, 32), to_signed(-687204285, 32), to_signed(-687362470, 32),
     to_signed(-687520629, 32), to_signed(-687678763, 32), to_signed(-687836872, 32), to_signed(-687994955, 32),
     to_signed(-688153013, 32), to_signed(-688311046, 32), to_signed(-688469054, 32), to_signed(-688627036, 32),
     to_signed(-688784993, 32), to_signed(-688942924, 32), to_signed(-689100831, 32), to_signed(-689258712, 32),
     to_signed(-689416567, 32), to_signed(-689574397, 32), to_signed(-689732202, 32), to_signed(-689889982, 32),
     to_signed(-690047736, 32), to_signed(-690205465, 32), to_signed(-690363168, 32), to_signed(-690520846, 32),
     to_signed(-690678499, 32), to_signed(-690836126, 32), to_signed(-690993728, 32), to_signed(-691151304, 32),
     to_signed(-691308855, 32), to_signed(-691466381, 32), to_signed(-691623881, 32), to_signed(-691781356, 32),
     to_signed(-691938805, 32), to_signed(-692096229, 32), to_signed(-692253627, 32), to_signed(-692411000, 32),
     to_signed(-692568348, 32), to_signed(-692725670, 32), to_signed(-692882966, 32), to_signed(-693040238, 32),
     to_signed(-693197483, 32), to_signed(-693354703, 32), to_signed(-693511898, 32), to_signed(-693669067, 32),
     to_signed(-693826211, 32), to_signed(-693983329, 32), to_signed(-694140422, 32), to_signed(-694297489, 32),
     to_signed(-694454530, 32), to_signed(-694611546, 32), to_signed(-694768537, 32), to_signed(-694925502, 32),
     to_signed(-695082441, 32), to_signed(-695239355, 32), to_signed(-695396243, 32), to_signed(-695553106, 32),
     to_signed(-695709943, 32), to_signed(-695866755, 32), to_signed(-696023541, 32), to_signed(-696180301, 32),
     to_signed(-696337036, 32), to_signed(-696493745, 32), to_signed(-696650429, 32), to_signed(-696807087, 32),
     to_signed(-696963719, 32), to_signed(-697120326, 32), to_signed(-697276907, 32), to_signed(-697433462, 32),
     to_signed(-697589992, 32), to_signed(-697746496, 32), to_signed(-697902975, 32), to_signed(-698059428, 32),
     to_signed(-698215855, 32), to_signed(-698372256, 32), to_signed(-698528632, 32), to_signed(-698684982, 32),
     to_signed(-698841307, 32), to_signed(-698997605, 32), to_signed(-699153879, 32), to_signed(-699310126, 32),
     to_signed(-699466348, 32), to_signed(-699622543, 32), to_signed(-699778714, 32), to_signed(-699934858, 32),
     to_signed(-700090977, 32), to_signed(-700247070, 32), to_signed(-700403137, 32), to_signed(-700559179, 32),
     to_signed(-700715194, 32), to_signed(-700871184, 32), to_signed(-701027149, 32), to_signed(-701183087, 32),
     to_signed(-701339000, 32), to_signed(-701494887, 32), to_signed(-701650748, 32), to_signed(-701806583, 32),
     to_signed(-701962393, 32), to_signed(-702118176, 32), to_signed(-702273934, 32), to_signed(-702429666, 32),
     to_signed(-702585372, 32), to_signed(-702741053, 32), to_signed(-702896707, 32), to_signed(-703052336, 32),
     to_signed(-703207939, 32), to_signed(-703363516, 32), to_signed(-703519067, 32), to_signed(-703674592, 32),
     to_signed(-703830092, 32), to_signed(-703985565, 32), to_signed(-704141013, 32), to_signed(-704296435, 32),
     to_signed(-704451830, 32), to_signed(-704607200, 32), to_signed(-704762544, 32), to_signed(-704917862, 32),
     to_signed(-705073155, 32), to_signed(-705228421, 32), to_signed(-705383661, 32), to_signed(-705538876, 32),
     to_signed(-705694064, 32), to_signed(-705849227, 32), to_signed(-706004363, 32), to_signed(-706159474, 32),
     to_signed(-706314559, 32), to_signed(-706469617, 32), to_signed(-706624650, 32), to_signed(-706779657, 32),
     to_signed(-706934638, 32), to_signed(-707089592, 32), to_signed(-707244521, 32), to_signed(-707399424, 32),
     to_signed(-707554301, 32), to_signed(-707709151, 32), to_signed(-707863976, 32), to_signed(-708018775, 32),
     to_signed(-708173547, 32), to_signed(-708328294, 32), to_signed(-708483015, 32), to_signed(-708637709, 32),
     to_signed(-708792378, 32), to_signed(-708947020, 32), to_signed(-709101636, 32), to_signed(-709256227, 32),
     to_signed(-709410791, 32), to_signed(-709565329, 32), to_signed(-709719841, 32), to_signed(-709874327, 32),
     to_signed(-710028787, 32), to_signed(-710183221, 32), to_signed(-710337628, 32), to_signed(-710492010, 32),
     to_signed(-710646365, 32), to_signed(-710800694, 32), to_signed(-710954997, 32), to_signed(-711109274, 32),
     to_signed(-711263525, 32), to_signed(-711417750, 32), to_signed(-711571948, 32), to_signed(-711726121, 32),
     to_signed(-711880267, 32), to_signed(-712034387, 32), to_signed(-712188481, 32), to_signed(-712342549, 32),
     to_signed(-712496590, 32), to_signed(-712650605, 32), to_signed(-712804594, 32), to_signed(-712958557, 32),
     to_signed(-713112494, 32), to_signed(-713266404, 32), to_signed(-713420288, 32), to_signed(-713574146, 32),
     to_signed(-713727978, 32), to_signed(-713881784, 32), to_signed(-714035563, 32), to_signed(-714189316, 32),
     to_signed(-714343043, 32), to_signed(-714496743, 32), to_signed(-714650417, 32), to_signed(-714804065, 32),
     to_signed(-714957687, 32), to_signed(-715111282, 32), to_signed(-715264851, 32), to_signed(-715418394, 32),
     to_signed(-715571910, 32), to_signed(-715725401, 32), to_signed(-715878864, 32), to_signed(-716032302, 32),
     to_signed(-716185713, 32), to_signed(-716339098, 32), to_signed(-716492457, 32), to_signed(-716645789, 32),
     to_signed(-716799095, 32), to_signed(-716952374, 32), to_signed(-717105627, 32), to_signed(-717258854, 32),
     to_signed(-717412054, 32), to_signed(-717565228, 32), to_signed(-717718376, 32), to_signed(-717871497, 32),
     to_signed(-718024592, 32), to_signed(-718177660, 32), to_signed(-718330702, 32), to_signed(-718483718, 32),
     to_signed(-718636707, 32), to_signed(-718789670, 32), to_signed(-718942606, 32), to_signed(-719095516, 32),
     to_signed(-719248400, 32), to_signed(-719401257, 32), to_signed(-719554087, 32), to_signed(-719706891, 32),
     to_signed(-719859669, 32), to_signed(-720012420, 32), to_signed(-720165145, 32), to_signed(-720317843, 32),
     to_signed(-720470515, 32), to_signed(-720623160, 32), to_signed(-720775779, 32), to_signed(-720928371, 32),
     to_signed(-721080937, 32), to_signed(-721233476, 32), to_signed(-721385989, 32), to_signed(-721538475, 32),
     to_signed(-721690935, 32), to_signed(-721843368, 32), to_signed(-721995775, 32), to_signed(-722148155, 32),
     to_signed(-722300508, 32), to_signed(-722452835, 32), to_signed(-722605136, 32), to_signed(-722757410, 32),
     to_signed(-722909657, 32), to_signed(-723061877, 32), to_signed(-723214072, 32), to_signed(-723366239, 32),
     to_signed(-723518380, 32), to_signed(-723670494, 32), to_signed(-723822582, 32), to_signed(-723974643, 32),
     to_signed(-724126677, 32), to_signed(-724278685, 32), to_signed(-724430667, 32), to_signed(-724582621, 32),
     to_signed(-724734549, 32), to_signed(-724886450, 32), to_signed(-725038325, 32), to_signed(-725190173, 32),
     to_signed(-725341994, 32), to_signed(-725493789, 32), to_signed(-725645557, 32), to_signed(-725797298, 32),
     to_signed(-725949013, 32), to_signed(-726100701, 32), to_signed(-726252362, 32), to_signed(-726403996, 32),
     to_signed(-726555604, 32), to_signed(-726707185, 32), to_signed(-726858740, 32), to_signed(-727010267, 32),
     to_signed(-727161768, 32), to_signed(-727313242, 32), to_signed(-727464690, 32), to_signed(-727616111, 32),
     to_signed(-727767504, 32), to_signed(-727918872, 32), to_signed(-728070212, 32), to_signed(-728221526, 32),
     to_signed(-728372813, 32), to_signed(-728524073, 32), to_signed(-728675306, 32), to_signed(-728826513, 32),
     to_signed(-728977692, 32), to_signed(-729128845, 32), to_signed(-729279971, 32), to_signed(-729431071, 32),
     to_signed(-729582143, 32), to_signed(-729733189, 32), to_signed(-729884208, 32), to_signed(-730035200, 32),
     to_signed(-730186165, 32), to_signed(-730337103, 32), to_signed(-730488014, 32), to_signed(-730638899, 32),
     to_signed(-730789757, 32), to_signed(-730940588, 32), to_signed(-731091392, 32), to_signed(-731242169, 32),
     to_signed(-731392919, 32), to_signed(-731543642, 32), to_signed(-731694339, 32), to_signed(-731845008, 32),
     to_signed(-731995651, 32), to_signed(-732146267, 32), to_signed(-732296855, 32), to_signed(-732447417, 32),
     to_signed(-732597952, 32), to_signed(-732748460, 32), to_signed(-732898941, 32), to_signed(-733049395, 32),
     to_signed(-733199822, 32), to_signed(-733350223, 32), to_signed(-733500596, 32), to_signed(-733650942, 32),
     to_signed(-733801261, 32), to_signed(-733951554, 32), to_signed(-734101819, 32), to_signed(-734252057, 32),
     to_signed(-734402269, 32), to_signed(-734552453, 32), to_signed(-734702610, 32), to_signed(-734852741, 32),
     to_signed(-735002844, 32), to_signed(-735152920, 32), to_signed(-735302970, 32), to_signed(-735452992, 32),
     to_signed(-735602987, 32), to_signed(-735752955, 32), to_signed(-735902896, 32), to_signed(-736052810, 32),
     to_signed(-736202697, 32), to_signed(-736352557, 32), to_signed(-736502390, 32), to_signed(-736652196, 32),
     to_signed(-736801974, 32), to_signed(-736951726, 32), to_signed(-737101450, 32), to_signed(-737251148, 32),
     to_signed(-737400818, 32), to_signed(-737550461, 32), to_signed(-737700077, 32), to_signed(-737849666, 32),
     to_signed(-737999228, 32), to_signed(-738148762, 32), to_signed(-738298270, 32), to_signed(-738447750, 32),
     to_signed(-738597203, 32), to_signed(-738746630, 32), to_signed(-738896028, 32), to_signed(-739045400, 32),
     to_signed(-739194745, 32), to_signed(-739344062, 32), to_signed(-739493352, 32), to_signed(-739642615, 32),
     to_signed(-739791851, 32), to_signed(-739941060, 32), to_signed(-740090241, 32), to_signed(-740239395, 32),
     to_signed(-740388522, 32), to_signed(-740537622, 32), to_signed(-740686694, 32), to_signed(-740835740, 32),
     to_signed(-740984758, 32), to_signed(-741133749, 32), to_signed(-741282712, 32), to_signed(-741431649, 32),
     to_signed(-741580558, 32), to_signed(-741729439, 32), to_signed(-741878294, 32), to_signed(-742027121, 32),
     to_signed(-742175921, 32), to_signed(-742324694, 32), to_signed(-742473439, 32), to_signed(-742622157, 32),
     to_signed(-742770848, 32), to_signed(-742919511, 32), to_signed(-743068147, 32), to_signed(-743216756, 32),
     to_signed(-743365338, 32), to_signed(-743513892, 32), to_signed(-743662419, 32), to_signed(-743810918, 32),
     to_signed(-743959390, 32), to_signed(-744107835, 32), to_signed(-744256253, 32), to_signed(-744404643, 32),
     to_signed(-744553005, 32), to_signed(-744701341, 32), to_signed(-744849649, 32), to_signed(-744997929, 32),
     to_signed(-745146182, 32), to_signed(-745294408, 32), to_signed(-745442606, 32), to_signed(-745590777, 32),
     to_signed(-745738921, 32), to_signed(-745887037, 32), to_signed(-746035126, 32), to_signed(-746183187, 32),
     to_signed(-746331221, 32), to_signed(-746479227, 32), to_signed(-746627206, 32), to_signed(-746775158, 32),
     to_signed(-746923082, 32), to_signed(-747070978, 32), to_signed(-747218847, 32), to_signed(-747366689, 32),
     to_signed(-747514503, 32), to_signed(-747662290, 32), to_signed(-747810049, 32), to_signed(-747957781, 32),
     to_signed(-748105485, 32), to_signed(-748253161, 32), to_signed(-748400811, 32), to_signed(-748548432, 32),
     to_signed(-748696026, 32), to_signed(-748843593, 32), to_signed(-748991132, 32), to_signed(-749138644, 32),
     to_signed(-749286127, 32), to_signed(-749433584, 32), to_signed(-749581013, 32), to_signed(-749728414, 32),
     to_signed(-749875788, 32), to_signed(-750023134, 32), to_signed(-750170453, 32), to_signed(-750317744, 32),
     to_signed(-750465007, 32), to_signed(-750612243, 32), to_signed(-750759451, 32), to_signed(-750906632, 32),
     to_signed(-751053785, 32), to_signed(-751200910, 32), to_signed(-751348008, 32), to_signed(-751495078, 32),
     to_signed(-751642121, 32), to_signed(-751789136, 32), to_signed(-751936123, 32), to_signed(-752083083, 32),
     to_signed(-752230015, 32), to_signed(-752376919, 32), to_signed(-752523796, 32), to_signed(-752670645, 32),
     to_signed(-752817466, 32), to_signed(-752964260, 32), to_signed(-753111025, 32), to_signed(-753257764, 32),
     to_signed(-753404474, 32), to_signed(-753551157, 32), to_signed(-753697812, 32), to_signed(-753844440, 32),
     to_signed(-753991040, 32), to_signed(-754137612, 32), to_signed(-754284156, 32), to_signed(-754430672, 32),
     to_signed(-754577161, 32), to_signed(-754723622, 32), to_signed(-754870056, 32), to_signed(-755016461, 32),
     to_signed(-755162839, 32), to_signed(-755309189, 32), to_signed(-755455511, 32), to_signed(-755601806, 32),
     to_signed(-755748072, 32), to_signed(-755894311, 32), to_signed(-756040522, 32), to_signed(-756186706, 32),
     to_signed(-756332861, 32), to_signed(-756478989, 32), to_signed(-756625089, 32), to_signed(-756771161, 32),
     to_signed(-756917205, 32), to_signed(-757063222, 32), to_signed(-757209210, 32), to_signed(-757355171, 32),
     to_signed(-757501104, 32), to_signed(-757647009, 32), to_signed(-757792886, 32), to_signed(-757938736, 32),
     to_signed(-758084557, 32), to_signed(-758230351, 32), to_signed(-758376116, 32), to_signed(-758521854, 32),
     to_signed(-758667564, 32), to_signed(-758813246, 32), to_signed(-758958900, 32), to_signed(-759104527, 32));  -- sfix32 [4096]

  -- Functions
  -- HDLCODER_TO_STDLOGIC 
  FUNCTION hdlcoder_to_stdlogic(arg: boolean) RETURN std_logic IS
  BEGIN
    IF arg THEN
      RETURN '1';
    ELSE
      RETURN '0';
    END IF;
  END FUNCTION;


  -- Signals
  SIGNAL stage_unsigned                   : unsigned(3 DOWNTO 0);  -- ufix4
  SIGNAL minResRX2FFTTwdlMapping_baseAddr : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL minResRX2FFTTwdlMapping_cnt      : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL minResRX2FFTTwdlMapping_octantReg1 : unsigned(2 DOWNTO 0);  -- ufix3
  SIGNAL minResRX2FFTTwdlMapping_twdlAddr_raw : unsigned(14 DOWNTO 0);  -- ufix15
  SIGNAL minResRX2FFTTwdlMapping_twdlAddrMap : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL minResRX2FFTTwdlMapping_twdl45Reg : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_dvldReg1 : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_dvldReg2 : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_maxCnt   : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL minResRX2FFTTwdlMapping_baseAddr_next : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL minResRX2FFTTwdlMapping_cnt_next : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL minResRX2FFTTwdlMapping_octantReg1_next : unsigned(2 DOWNTO 0);  -- ufix3
  SIGNAL minResRX2FFTTwdlMapping_twdlAddr_raw_next : unsigned(14 DOWNTO 0);  -- ufix15
  SIGNAL minResRX2FFTTwdlMapping_twdlAddrMap_next : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL minResRX2FFTTwdlMapping_twdl45Reg_next : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_dvldReg1_next : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_dvldReg2_next : std_logic;
  SIGNAL minResRX2FFTTwdlMapping_maxCnt_next : unsigned(13 DOWNTO 0);  -- ufix14
  SIGNAL twdlAddr                         : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL twdlAddrVld                      : std_logic;
  SIGNAL twdlOctant                       : unsigned(2 DOWNTO 0);  -- ufix3
  SIGNAL twdl45                           : std_logic;
  SIGNAL twiddleS_re                      : signed(31 DOWNTO 0);  -- sfix32_En30
  SIGNAL twiddleReg_re                    : signed(31 DOWNTO 0);  -- sfix32_En30
  SIGNAL twiddleS_im                      : signed(31 DOWNTO 0);  -- sfix32_En30
  SIGNAL twiddleReg_im                    : signed(31 DOWNTO 0);  -- sfix32_En30
  SIGNAL twdlOctantReg                    : unsigned(2 DOWNTO 0);  -- ufix3
  SIGNAL twdl45Reg                        : std_logic;
  SIGNAL twdl_re_tmp                      : signed(31 DOWNTO 0);  -- sfix32_En30
  SIGNAL twdl_im_tmp                      : signed(31 DOWNTO 0);  -- sfix32_En30

BEGIN
  stage_unsigned <= unsigned(stage);

  -- minResRX2FFTTwdlMapping
  minResRX2FFTTwdlMapping_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      minResRX2FFTTwdlMapping_octantReg1 <= to_unsigned(16#0#, 3);
      minResRX2FFTTwdlMapping_twdlAddr_raw <= to_unsigned(16#0000#, 15);
      minResRX2FFTTwdlMapping_twdlAddrMap <= to_unsigned(16#000#, 12);
      minResRX2FFTTwdlMapping_twdl45Reg <= '0';
      minResRX2FFTTwdlMapping_dvldReg1 <= '0';
      minResRX2FFTTwdlMapping_dvldReg2 <= '0';
      minResRX2FFTTwdlMapping_baseAddr <= to_unsigned(16#0000#, 14);
      minResRX2FFTTwdlMapping_cnt <= to_unsigned(16#3FFF#, 14);
      minResRX2FFTTwdlMapping_maxCnt <= to_unsigned(16#0000#, 14);
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        IF syncReset = '1' THEN
          minResRX2FFTTwdlMapping_octantReg1 <= to_unsigned(16#0#, 3);
          minResRX2FFTTwdlMapping_twdlAddr_raw <= to_unsigned(16#0000#, 15);
          minResRX2FFTTwdlMapping_twdlAddrMap <= to_unsigned(16#000#, 12);
          minResRX2FFTTwdlMapping_twdl45Reg <= '0';
          minResRX2FFTTwdlMapping_dvldReg1 <= '0';
          minResRX2FFTTwdlMapping_dvldReg2 <= '0';
          minResRX2FFTTwdlMapping_baseAddr <= to_unsigned(16#0000#, 14);
          minResRX2FFTTwdlMapping_cnt <= to_unsigned(16#3FFF#, 14);
          minResRX2FFTTwdlMapping_maxCnt <= to_unsigned(16#0000#, 14);
        ELSE 
          minResRX2FFTTwdlMapping_baseAddr <= minResRX2FFTTwdlMapping_baseAddr_next;
          minResRX2FFTTwdlMapping_cnt <= minResRX2FFTTwdlMapping_cnt_next;
          minResRX2FFTTwdlMapping_octantReg1 <= minResRX2FFTTwdlMapping_octantReg1_next;
          minResRX2FFTTwdlMapping_twdlAddr_raw <= minResRX2FFTTwdlMapping_twdlAddr_raw_next;
          minResRX2FFTTwdlMapping_twdlAddrMap <= minResRX2FFTTwdlMapping_twdlAddrMap_next;
          minResRX2FFTTwdlMapping_twdl45Reg <= minResRX2FFTTwdlMapping_twdl45Reg_next;
          minResRX2FFTTwdlMapping_dvldReg1 <= minResRX2FFTTwdlMapping_dvldReg1_next;
          minResRX2FFTTwdlMapping_dvldReg2 <= minResRX2FFTTwdlMapping_dvldReg2_next;
          minResRX2FFTTwdlMapping_maxCnt <= minResRX2FFTTwdlMapping_maxCnt_next;
        END IF;
      END IF;
    END IF;
  END PROCESS minResRX2FFTTwdlMapping_process;

  minResRX2FFTTwdlMapping_output : PROCESS (dMemOutDly_vld, initIC, minResRX2FFTTwdlMapping_baseAddr,
       minResRX2FFTTwdlMapping_cnt, minResRX2FFTTwdlMapping_dvldReg1,
       minResRX2FFTTwdlMapping_dvldReg2, minResRX2FFTTwdlMapping_maxCnt,
       minResRX2FFTTwdlMapping_octantReg1, minResRX2FFTTwdlMapping_twdl45Reg,
       minResRX2FFTTwdlMapping_twdlAddrMap,
       minResRX2FFTTwdlMapping_twdlAddr_raw, stage_unsigned)
    VARIABLE octant : unsigned(2 DOWNTO 0);
    VARIABLE sub_cast : signed(31 DOWNTO 0);
    VARIABLE sub_temp : signed(31 DOWNTO 0);
    VARIABLE sub_cast_0 : signed(16 DOWNTO 0);
    VARIABLE sub_temp_0 : signed(16 DOWNTO 0);
    VARIABLE sub_cast_1 : signed(16 DOWNTO 0);
    VARIABLE sub_temp_1 : signed(16 DOWNTO 0);
    VARIABLE sub_cast_2 : signed(31 DOWNTO 0);
    VARIABLE sub_temp_2 : signed(31 DOWNTO 0);
    VARIABLE sub_cast_3 : signed(31 DOWNTO 0);
    VARIABLE sub_temp_3 : signed(31 DOWNTO 0);
  BEGIN
    sub_temp := to_signed(0, 32);
    sub_temp_0 := to_signed(16#00000#, 17);
    sub_temp_1 := to_signed(16#00000#, 17);
    sub_temp_2 := to_signed(0, 32);
    sub_temp_3 := to_signed(0, 32);
    sub_cast := to_signed(0, 32);
    sub_cast_0 := to_signed(16#00000#, 17);
    sub_cast_1 := to_signed(16#00000#, 17);
    sub_cast_2 := to_signed(0, 32);
    sub_cast_3 := to_signed(0, 32);
    minResRX2FFTTwdlMapping_baseAddr_next <= minResRX2FFTTwdlMapping_baseAddr;
    minResRX2FFTTwdlMapping_cnt_next <= minResRX2FFTTwdlMapping_cnt;
    minResRX2FFTTwdlMapping_twdlAddrMap_next <= minResRX2FFTTwdlMapping_twdlAddrMap;
    minResRX2FFTTwdlMapping_twdl45Reg_next <= minResRX2FFTTwdlMapping_twdl45Reg;
    minResRX2FFTTwdlMapping_maxCnt_next <= minResRX2FFTTwdlMapping_maxCnt;
    minResRX2FFTTwdlMapping_dvldReg2_next <= minResRX2FFTTwdlMapping_dvldReg1;
    minResRX2FFTTwdlMapping_dvldReg1_next <= dMemOutDly_vld;
    CASE minResRX2FFTTwdlMapping_twdlAddr_raw IS
      WHEN "001000000000000" =>
        octant := to_unsigned(16#0#, 3);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '1';
      WHEN "010000000000000" =>
        octant := to_unsigned(16#1#, 3);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '0';
      WHEN "011000000000000" =>
        octant := to_unsigned(16#2#, 3);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '1';
      WHEN "100000000000000" =>
        octant := to_unsigned(16#3#, 3);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '0';
      WHEN "101000000000000" =>
        octant := to_unsigned(16#4#, 3);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '1';
      WHEN OTHERS => 
        octant := minResRX2FFTTwdlMapping_twdlAddr_raw(14 DOWNTO 12);
        minResRX2FFTTwdlMapping_twdl45Reg_next <= '0';
    END CASE;
    minResRX2FFTTwdlMapping_octantReg1_next <= octant;
    CASE octant IS
      WHEN "000" =>
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= minResRX2FFTTwdlMapping_twdlAddr_raw(11 DOWNTO 0);
      WHEN "001" =>
        sub_cast_0 := signed(resize(minResRX2FFTTwdlMapping_twdlAddr_raw, 17));
        sub_temp_0 := to_signed(16#02000#, 17) - sub_cast_0;
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= unsigned(sub_temp_0(11 DOWNTO 0));
      WHEN "010" =>
        sub_cast_1 := signed(resize(minResRX2FFTTwdlMapping_twdlAddr_raw, 17));
        sub_temp_1 := sub_cast_1 - to_signed(16#02000#, 17);
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= unsigned(sub_temp_1(11 DOWNTO 0));
      WHEN "011" =>
        sub_cast_2 := signed(resize(minResRX2FFTTwdlMapping_twdlAddr_raw & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0', 32));
        sub_temp_2 := to_signed(67108864, 32) - sub_cast_2;
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= unsigned(sub_temp_2(23 DOWNTO 12));
      WHEN "100" =>
        sub_cast_3 := signed(resize(minResRX2FFTTwdlMapping_twdlAddr_raw & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0', 32));
        sub_temp_3 := sub_cast_3 - to_signed(67108864, 32);
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= unsigned(sub_temp_3(23 DOWNTO 12));
      WHEN OTHERS => 
        sub_cast := signed(resize(minResRX2FFTTwdlMapping_twdlAddr_raw & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0', 32));
        sub_temp := to_signed(100663296, 32) - sub_cast;
        minResRX2FFTTwdlMapping_twdlAddrMap_next <= unsigned(sub_temp(23 DOWNTO 12));
    END CASE;
    minResRX2FFTTwdlMapping_twdlAddr_raw_next <= resize(unsigned'(minResRX2FFTTwdlMapping_baseAddr(0) & minResRX2FFTTwdlMapping_baseAddr(1) & minResRX2FFTTwdlMapping_baseAddr(2) & minResRX2FFTTwdlMapping_baseAddr(3) & minResRX2FFTTwdlMapping_baseAddr(4) & minResRX2FFTTwdlMapping_baseAddr(5) & minResRX2FFTTwdlMapping_baseAddr(6) & minResRX2FFTTwdlMapping_baseAddr(7) & minResRX2FFTTwdlMapping_baseAddr(8) & minResRX2FFTTwdlMapping_baseAddr(9) & minResRX2FFTTwdlMapping_baseAddr(10) & minResRX2FFTTwdlMapping_baseAddr(11) & minResRX2FFTTwdlMapping_baseAddr(12) & minResRX2FFTTwdlMapping_baseAddr(13)), 15);
    IF ( NOT initIC) = '1' THEN 
      IF (dMemOutDly_vld AND hdlcoder_to_stdlogic(minResRX2FFTTwdlMapping_cnt = to_unsigned(16#0000#, 14))) = '1' THEN 
        minResRX2FFTTwdlMapping_baseAddr_next <= minResRX2FFTTwdlMapping_baseAddr + to_unsigned(16#0001#, 14);
      END IF;
    ELSE 
      minResRX2FFTTwdlMapping_baseAddr_next <= to_unsigned(16#0000#, 14);
    END IF;
    IF ( NOT initIC) = '1' THEN 
      IF dMemOutDly_vld = '1' THEN 
        IF minResRX2FFTTwdlMapping_cnt = to_unsigned(16#0000#, 14) THEN 
          minResRX2FFTTwdlMapping_cnt_next <= minResRX2FFTTwdlMapping_maxCnt;
        ELSE 
          minResRX2FFTTwdlMapping_cnt_next <= minResRX2FFTTwdlMapping_cnt - to_unsigned(16#0001#, 14);
        END IF;
      END IF;
    ELSIF stage_unsigned = to_unsigned(16#0#, 4) THEN 
      minResRX2FFTTwdlMapping_maxCnt_next <= to_unsigned(16#3FFF#, 14);
      minResRX2FFTTwdlMapping_cnt_next <= to_unsigned(16#3FFF#, 14);
    ELSE 
      minResRX2FFTTwdlMapping_cnt_next <= minResRX2FFTTwdlMapping_maxCnt srl 1;
      minResRX2FFTTwdlMapping_maxCnt_next <= minResRX2FFTTwdlMapping_maxCnt srl 1;
    END IF;
    twdlAddr <= minResRX2FFTTwdlMapping_twdlAddrMap;
    twdlAddrVld <= minResRX2FFTTwdlMapping_dvldReg2;
    twdlOctant <= minResRX2FFTTwdlMapping_octantReg1;
    twdl45 <= minResRX2FFTTwdlMapping_twdl45Reg;
  END PROCESS minResRX2FFTTwdlMapping_output;


  -- Twiddle ROM1
  twiddleS_re <= Twiddle_re_table_data(to_integer(twdlAddr));

  TWIDDLEROM_RE_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      twiddleReg_re <= to_signed(0, 32);
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        twiddleReg_re <= twiddleS_re;
      END IF;
    END IF;
  END PROCESS TWIDDLEROM_RE_process;


  -- Twiddle ROM2
  twiddleS_im <= Twiddle_im_table_data(to_integer(twdlAddr));

  TWIDDLEROM_IM_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      twiddleReg_im <= to_signed(0, 32);
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        twiddleReg_im <= twiddleS_im;
      END IF;
    END IF;
  END PROCESS TWIDDLEROM_IM_process;


  intdelay_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      twdlOctantReg <= to_unsigned(16#0#, 3);
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        IF syncReset = '1' THEN
          twdlOctantReg <= to_unsigned(16#0#, 3);
        ELSE 
          twdlOctantReg <= twdlOctant;
        END IF;
      END IF;
    END IF;
  END PROCESS intdelay_process;


  intdelay_1_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      twdl45Reg <= '0';
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        IF syncReset = '1' THEN
          twdl45Reg <= '0';
        ELSE 
          twdl45Reg <= twdl45;
        END IF;
      END IF;
    END IF;
  END PROCESS intdelay_1_process;


  -- Radix22TwdlOctCorr
  Radix22TwdlOctCorr_output : PROCESS (twdl45Reg, twdlOctantReg, twiddleReg_im, twiddleReg_re)
    VARIABLE twdlIn_re : signed(31 DOWNTO 0);
    VARIABLE twdlIn_im : signed(31 DOWNTO 0);
    VARIABLE cast : signed(32 DOWNTO 0);
    VARIABLE cast_0 : signed(32 DOWNTO 0);
    VARIABLE cast_1 : signed(32 DOWNTO 0);
    VARIABLE cast_2 : signed(32 DOWNTO 0);
    VARIABLE cast_3 : signed(32 DOWNTO 0);
    VARIABLE cast_4 : signed(32 DOWNTO 0);
    VARIABLE cast_5 : signed(32 DOWNTO 0);
    VARIABLE cast_6 : signed(32 DOWNTO 0);
    VARIABLE cast_7 : signed(32 DOWNTO 0);
    VARIABLE cast_8 : signed(32 DOWNTO 0);
    VARIABLE cast_9 : signed(32 DOWNTO 0);
    VARIABLE cast_10 : signed(32 DOWNTO 0);
  BEGIN
    cast_0 := to_signed(0, 33);
    cast_2 := to_signed(0, 33);
    cast_4 := to_signed(0, 33);
    cast_6 := to_signed(0, 33);
    cast_8 := to_signed(0, 33);
    cast_10 := to_signed(0, 33);
    cast := to_signed(0, 33);
    cast_1 := to_signed(0, 33);
    cast_3 := to_signed(0, 33);
    cast_5 := to_signed(0, 33);
    cast_7 := to_signed(0, 33);
    cast_9 := to_signed(0, 33);
    twdlIn_re := twiddleReg_re;
    twdlIn_im := twiddleReg_im;
    IF twdl45Reg = '1' THEN 
      CASE twdlOctantReg IS
        WHEN "000" =>
          twdlIn_re := to_signed(759250125, 32);
          twdlIn_im := to_signed(-759250125, 32);
        WHEN "010" =>
          twdlIn_re := to_signed(-759250125, 32);
          twdlIn_im := to_signed(-759250125, 32);
        WHEN "100" =>
          twdlIn_re := to_signed(-759250125, 32);
          twdlIn_im := to_signed(759250125, 32);
        WHEN OTHERS => 
          twdlIn_re := to_signed(759250125, 32);
          twdlIn_im := to_signed(-759250125, 32);
      END CASE;
    ELSE 
      CASE twdlOctantReg IS
        WHEN "000" =>
          NULL;
        WHEN "001" =>
          cast := resize(twiddleReg_im, 33);
          cast_0 :=  - (cast);
          twdlIn_re := cast_0(31 DOWNTO 0);
          cast_5 := resize(twiddleReg_re, 33);
          cast_6 :=  - (cast_5);
          twdlIn_im := cast_6(31 DOWNTO 0);
        WHEN "010" =>
          twdlIn_re := twiddleReg_im;
          cast_7 := resize(twiddleReg_re, 33);
          cast_8 :=  - (cast_7);
          twdlIn_im := cast_8(31 DOWNTO 0);
        WHEN "011" =>
          cast_1 := resize(twiddleReg_re, 33);
          cast_2 :=  - (cast_1);
          twdlIn_re := cast_2(31 DOWNTO 0);
          twdlIn_im := twiddleReg_im;
        WHEN "100" =>
          cast_3 := resize(twiddleReg_re, 33);
          cast_4 :=  - (cast_3);
          twdlIn_re := cast_4(31 DOWNTO 0);
          cast_9 := resize(twiddleReg_im, 33);
          cast_10 :=  - (cast_9);
          twdlIn_im := cast_10(31 DOWNTO 0);
        WHEN OTHERS => 
          twdlIn_re := twiddleReg_im;
          twdlIn_im := twiddleReg_re;
      END CASE;
    END IF;
    twdl_re_tmp <= twdlIn_re;
    twdl_im_tmp <= twdlIn_im;
  END PROCESS Radix22TwdlOctCorr_output;


  twdl_re <= std_logic_vector(twdl_re_tmp);

  twdl_im <= std_logic_vector(twdl_im_tmp);

END rtl;

